��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t�������.NT��8\�Q��ȍ�������H�V�&�bO�t0ķ��~?�c��d�]L}�L�`������������	��f���|cl����B��x�E.�		��@2��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HCZ�C�Ru�����[H��22P^��{������6�a�WN8�L�u�E�>F5��o{�R~�Y\m�Ȕ.��K�Q�ց2.����/8��cG��B�+�%Y栠��'ޭ�--j��7��ml.���~j�n����©�kh�ؐ��=?�^J.W�Ս�8�"n�B,�U��,�qQ�0��'vI�?�֐`6^�fv����x�Bڻ�.8��9X\�7������TиEm�;����ME`���͎�ݱ�tĳ�U�����Qw�_� �6Тj�&[+�{˲
���Vŋ3`��9b�ϡ<|�9 L�p����\�%p�+aNߎ��l�;�0�)��Q�؍a5O<�8k�P��gM5�5�+}���?�h��ᤊ7d?4��_ڼ������E)�N˴vUK���Z1����)�?�APB�7���p����-DҨ���DV+Vy��3��R��T��E���sǊ�����j���JD#���!����C�Ʋ#�+H�6�8s��s]kFO_҈��r�b�L�* X�+Ƚ�b�V�P��E�2A��%�5n�	���l�#4\��B����?"ʕ����4@e�y��loa4#��z�hM��y(��3�贶�)�Mű� ��$G���I�f
)U�Khg�-4	)&I;�Ť�c ��!��n���?w�q�O#Y1�b9�x�bub�I�4Z��?E*T��9������#�W����#'��_�T=0>-G�{��j��U�O��8��5���J��t�/����=I��|��D3�T�4�$;8,��Ç�#Qk.QwdC���ш���MV�"�]�VW����)�W��f��FCL6�Y��15B~y#���Hv PZM��X#e;1�\LsɄ��F��n;��OM�Q�&<�i���9w��]�bw�O�`�o��~ZR�+TbuL~Ԇo��tht�β����"g��%�����z5�S����͡��:�����"�f� nH�$$7)O:^cS��(��g]�#35I-S(͋��u�/��pH#�vp�����X�#�@b?���r��I�[x���>'M�yL� |߯���:�rLZwI��c�R�ڥk
�yIC���!<��kx���ă��.Q��b1S�(�t��5�wtn�M��U�m8������1 U���,�x�0B3�b∊�Z��:��U�Z\��4Y���(�N���sQ�/��e�����%��Pkr5����c� R5�5l����y�a���mV��7nr�|/���/�]3?τ��#f�|_��WU��e\��٢!����Ԥ[�u��4}xk-"I��$ix�/Q.^d��\;d/%��9� �(�`�8�ҧ��� ��。䃙C�Cў�	L9�mU5Y8�t?����3fV<���A��(E]���BRZٙ��n("�����n�U�REw�U�@���U.��?�HVQ$�iǃiEr���V�[���2r��6~f*�����!�Iq����*�>�;�.���У�l���t�rˣ�W�4�z�������?�)����y?��'m���}wY2Ц���Ou�L��P�>���Et�2Q��9c\�e��9P���,��QD,ܬ�9�0C�ü2;?�)��[gg����[�	t���\BnZ�}cu�BŦ�AUDi$,=�B��p�0
?�X/���������Q�a6�"�#r鵃�֟?��Z"�mg��@���ِ�����me��X�朮�zܱIh�L6=S���HֈO�R�b��9���E:֝���V���7�$j41 �ٷS�2�w}��T]OrW�ۥV��T�{Ѷ_�X���D�-��f�Y��8�m�G߉�o�ڳɌ#O�E`$Lg���񮈺>��������c���kD ������cJ*tȔ�a����@���Ƅh+��@�%��oaxs��e�R5r*�~[�D/jRy�$V��� �G����W`x���<���y��H�����g C݄zZu6!�'��B#<��񧈝���c�un`�^�1�(2�����F��,�i�񈁛F�nYl�:�/�ۇ�����d)Rݔ ��\�?tnEq���55a:#A�a�xz=J⟐��d~�p��BO��r��<����
�c��lA�W�i�fgt·V���jN����2�u�ic����zX⒌0`��|���e��4�|���2i1�|�'e^*��t�g_��i�����a��4dIkl,E}�AQjM����w�+p�z�r�������ڦD��U�t+�|N���eW�.��϶+݀O�4�]M$T��nu�B�=_$��iGMSp Ѣ�T��r�*%ݘW�F��~����C�h�wt����W��c8�K�QNMd��>�]"��&��A0FkB��˒G�5�����0UP�1���.����
m�,���w�gt[�oB ���*����c��B���DT�C��~�/��𸇡� 1��XW�����k���m��;�euh�^�P�ձz�^�T�{k����1	@� ���D�{��/���-��lĨ��3QƠ�I5��R�˥OD�{��P���2�]e)�N�o�q�Sc\wi ���i���eL�񃨞C�Ր��qg�K��2U�x2l4g��NN��*���0u�x��1��ׄr�Z���.|_O�ڶHyE?��y�x	$*��I"����Q�х���Q��m����4��9s�Vxk����x�~�rN@���|i�k$W���w�����e0x��w�%�威 �BW��v5x�<(�a�j��4Ô��X�&L,(ы��90���*�˷���J�Vj�Z�sZ������:�"�c�S({	�=ʝ&��]H�߶X:.
��A��V��8���:ro)C��v�S�a� ]<��:7���2\���E[W�+��&9k��hCT�f�vmC�DX��`yUU�}�vd��(��\?^` �)�S�]y+�onN�35N�̋M>8�ոUt�21��r(��0����.��)?�j���
���)�(=OWʂ &m�\�-*m֮������D��tu������%+�)��S�l� 'fGrJ� ��}��b�l��S�h6;JZ��^���2�@�$*��5=�;ޜ���靜�-�������U�9�i.�,8m�^��(�C�"u�v�{>��t��|Q$b/
���=���l��\o��	MT��ER\Q������n@_Xs,�6]���� ��h��C�+*��"��oG��9 ���&��ן7�'�D7���Y�b�ֳ?�,�m1��x!�8gj�5�ϻ��b�oz�����
n)�!3���T��{�k?�+dcz�&O?�0(���sLQ�dfp��%ҧ1 ���Z?�V?�W��5��g]��)3�/��jH7l�-�_����N���i�S�ZVj�H�A}�|�dw����.ڻw���fK���=f�������".Oj"
��%��Y$x��9���`w��O��s�e��a��9`��k���S�~�g=B�SO=��(�0�P���J�8q�9����%rpƔ�8�;/-�Ʋ�s�9H������y
����N���x⭇��3�Y'���ʳډx�mpyB��ڙЯ��Z� ly?�y�Z�k@��cB��V������dJ:�w-ޞ��E)^��%��.{���sO%�cM��=���p�,��j�4��ȴU]"��${�I81��z�Q1�S,17��|���k���z�+���Uw���V���2��-����d�mȦ�\��>��܎���P��������t��L�X�c�(~�.J S_���i(V�0�V=a�i?��'��/yo�m2��Y�^ऻ��ȝ��[�@8���_��� 'ݭ�u����́��œ�ȑb�m��|3ǳ>�;|,��?vj�!�N�5���6�q��BX.&�rLa\J�X{����	�8 �\}S0-m欏i?�I�K��	���ɨ
�}s��H�`����g>p����Y4�9#'V��,���o�ˮ�~H �9�К� wBP��Э��p�Q�У{?�Cn�}�_D\E�ƅ瘍EӼ�m��2�e�ք�^ٯ"��V+[�C
�W"�@�F�9"�øV�A'�e�\��������oҍ��a�읢�K�я�l}����� $3^N#^k�j��ӊ�ߴv1[�;�ySt���a腇y�(�r�-6��K��U�O^��b�Ѡ���k�*��I�������0k�q����ʁ;��#k�I���3�]1��0#-3���{`AyE�t�P��S�>���c�.����+Slږ�~���W��$�Y,�H
�2�UO�a.NCw��*�Ѽ��$��9� հt0G���]/i�`[|\X�#)�4�`)���r�u$���5ֶ�z�)�+�3��lƥۊ�1�p���m�=T&Ι�A�"ضLzۤ�˗�[|�paU0�
Ů+ўb���#J��J0(F̎JG@��0�K��ގd!k$.3�$��w��n?]vf�;�R/�����!��ѷ��3@����Ϥ��p�\���E���>L?U?G�~ca�*��{k6�u�#1�����@h��Z;T(xD�0v ?dX�޾~4�!c��=�xX*���_A� GP�؇����������E[�Բ�]؍x`��߮2��=qr��ˤI^INc�/� Z�] ������OGwD���_5��v��&dfT$ (7� '*e��u�{h�o�4�p��<bC�A��Y�q�y����m#�fY94pz�K&�Y}Y�ufD5���1o�EN�;��1��qPF|�w ���G��;��w�y�}��.��I̥Lh��\�,���\�ǫ�%�ל{=X,6�'_����`ю�}�K�ݠ:ޘX=p������.�����?�!P����f��y��F��̤���u��_�x�I��t�Dx���<�� �)N�:�^|Y�蠱{�Lh���˰Z`�T"���ׄ/�� 6+�f�p�J2ϓ��;u(��aO]ˁ�������4��2�f�~���'�4������q4��x�{����,����LXP����m�hy�Wu.�J����1H�p7��8�X���M�jWf�����AYċ`�l,c�?� (�U�^���S�C�Qp�8�Ǵ&���ku��9���W�&����|�W��Q���&L}�N�_�pE��傁q	s������s�-Z�V.U��%U����k�R�л�4���\&��r�tI�����V�	3!u��rn;�@_�2��y|��`ȦL9n*q�[?�B���mM�Y�؎�T��~3�*L�AkxE��5V�6p��4g�ң��InJaX�G�sc^�w���Tc���)*��jal�F�w�W&k�EK~��}H)WC[tW����S�pO��O_��=#�����ђK�'��ܛn	���1�Ax˸��ɮW��!:G���s�e.���Ɍ�F�"5f���념�7�ZIbxj�tGuE���Mz7r�K��)�W(o��K������]��{��ءk+-���m���LZ�hg��޽9{@�� $�������q�v-����̣�n��ϝ7]�_=�mceL���0%�tw�ɵb-	fR�!���=,đx���f�}���u���Hl>Uo9��Q�gi��u��_���"�ʝ �O�
/�L��t*o�}�km�ʇ�!�yR�/7�fK������� ���	CZ��  x��'T5����mن:45lэI�;X�^T.v�	k1�~9/���������K�oՀ�XG"@|�D��n,,
��m���K���CzH�G��d'�.�-M��l+�d\[��צ��4t��Jz����<�T�GV��Nq0e��!U��*���w���m������G��)���X\���w�g;²
U�8�A��?~��{r������g�&qó̙D��ԅ�љ�:����\� 슶=��bX�(�pqv@{k���y�[��K� fj&å/�Cy0��`f�V9ә��2>l{0#ɶǋ���?&f�d�/�C�����KƇPL��1w��o���B�L3��^	�ܖ�����.Q-/�����s�b�]z�*���P,<��@oY^�R؈}��!��E[J4C~�	��X�M�W�>�1f��8�]���������jq���|�Â*������\
��7����`�J��T(�0yƿҊ��8�ؿ67j���֪1-������>��������[�JB�^;Rb~P�-��T|�ϔ�o���9�㏔n�G_т�^b����硙bLl�z������*�O�|�E���8aMsi^��;�z(����̿:a�K��e������fa�~H���Vu>�Ul7��ɮE�
��'Уç��[���[d�=�����kA�v�A�Ɩl������Vڢ�ze3/ܼ���%����(�iǌ�ie���?p��-��z�#���^��l��9#�BZ���y�c;�Rw;~1 �%����G������,ޑbHZ�,���"tb��[e��H��кmN;o�>x��a�������_~I&��&�Ӵ�C��n�A��-d�"}>ӊ�j��Rp6�',C�>�����|��>�9�={��A!w�a�ث.���uV@���#ʃ9*�8��2\F�`��dN����7#zeo��5ޟ��S�ɂX�XX�`���|7�b)�x�d��r1�@j�̜͌ �u�X�������9$�8p�Z����\�ު����T���ir���I��f0M&p���V�R�7\���<M7�ͤf���;�o�Nb���}�U�<����������kQ9�\��h̕$���v��U��`�u��ަ�ു��'y��uBh@�M�Wи[���b5��
�]_��) A����vC�PC�Fa�?_���t����������xu��Y�ˢ+����h��h�M��6�w}�%�����Db)8����zE���!.h��Z�d3v+~�
tBv����UJ�}�֢�$�~�n���8O��N[���:���q��) ��
�5嘍�����x��cu������{�чX��Kj^K<��/�	K2.x|������q7�}QK�i@�Q`����G}���|fē��n��l��h��㩿��&��F��z�%;
~�f��i���k��]����+]�)�0�<� b�	s+�!�1M�nө#߾:��V�5#������΅�
G�2�Վp����Jx�;ԍ�PiS^�;�`0Ƭ���k�� ��(�s��W���h�PyP�P\�c;fb�9�f�:�Z�z���#�g���f8�&|��Y݁�|h=���6�M��U�����W3H7���ܪd��Xll��O���	~!��I�/���#��1f�.e���7�)�L�O�z���Ρ��{��@��yT���h����)ӕf�K�?W�#J��$�L=1 �QGMt�yl�U_&"1�U�Mُ�C� ���OCa�c�:���,=�Hϧ�_v�f�wN��0��� ������\��ܔ0؄�@䴥��O�Ƌ��1���f;E{�SOScD�b8��k�u-�?y�UH �>N=�ځoXk��<FL���8S������`�5@��R��K��G�6/�Y���d�fb�l�t�MC@$�Q�XUw&�P��6h�DЫJɃ8>� Mp�����Q� j�~�0Z���$隐e�kĮ��~�A��H�M]Õ�Ft<Q��lr�1���-D�Y��m@ہ$���h�Hv�K�������X�i�
�r��w ˺B�����1^��j�dL�.����.kS���+fd�4x.���  GU���ů�������7<e�iZ��[�Jo�G�,��.n=��ư����j�pr�K�Ny��n,p�=��^Q���&����7��쎝6�J%�{��AVRZ��2�X��ia�޳	TD��K�Z n��+6-�7�
h티a|&�N�ر�9����v�����l�<b�JN$\/��,B�VT r7F<�j�[��|�����	��H(
�f$Y�ڦ)$X9O*a�d�8���x�BԢ��d<H\Ϝ�(nE�w� ���4��az�۶Z��J݊��p{��\����(cQ�,YT;�U}91O�\��Տ� d梳�!�df��)�W��/ ����-�������x	��7�p����S�X������#�����NL��g�������\c8�%'!�� ��e/��(�G���j
Cʰ�#��e�����<X���']�颧�h���9�g�`��͛�$L����D�����j��b�J�#2���Տ�������1�e�g(�@x��*��@o�.��B������7�Hi|6���X��s���^h��a�`S��-}��n����ͷЅeg!~�l?��=���	����g�Ǖ��}&@��P�-�|-�}�58��k�;7�Y�C�+�0������x��)�fC���+��as��W����D1Û����P��#"���m3���]�0`�g���T��>D�P`�n@z<
7_|�:��aI1���l[�J�]Y�A=0��x�=�,����&r��Trv�������9,d����>���f�E����|���#>َ���g���2i�'uE����W���3��s)?>�d�#�AE�HB���;�zq����T��k�G�s��#L��#ezޗ�������+^�f���q������	ډ&f���y=���X�f�}�H�((ۤ�|,9�GX8���ucwl@[Y0�:�l���
�0L ��_��n�
�N�Nē���@�p��s�C�b�?��R!��h#���d+#�)/�����"��|��{��""X��YX�F-b��{]﬛A���p�gF��E�1T��_9L���LG�ws��m�k�ǟ}͛e�!+�q���v��!�	�Y䨿�#ѷ߹����%ө�\W��8{��t�:��N_;�b�ֵ���*Gh'���6�?�]v�q�g�?ez�;6��>�W�0����0i��u
��{o��Vk�g�/l��/�����]tW�ɦ{}���-�cW�g �[ჲC�4F�6��蠣�����s��X%}�j}����K$9.�e�J�rmv�<G�c��T~�xL�@����ٜV�aI�,+f5))�0'Y�v/N�h7���ߜ�%Ӗ��3dz雌s��=���7 �vS�p}���, ����x�u�Jɼk��o_�Q�^Oq`܈'O���`9�q�:Ns��\���QO�^���:A�C�ϔb��+#�4�Q��}r^�v��G�Lz ��ŵ �f�*brb4�����5_�aXb���S�G䨤IpB��{c���HͣB�I�]� ��Q�q��Ô����6���Ta����Y���, �@���8��>��1�ؒ� �P{�]C��	r�\ORȐ�j�~��WCeJ�i�Nzß��j_qf.o�������xL��9�3p4�/���s���`�i�~]�:&�(��L�S\�7�pVD|D�����3klY���X�XC���\�ʍ���{�����m�g�Sc����/X�^�;L��3` [��ph�� ��Z<o�gܪ�po��2x��}��JA�d�"M�Q�1�H��Q����<Hc1�L#l�m߻�L@!�5[�8��L�$����#����V��E��2ϡ��Wn_��0f�[�E�$�_)fě�&Gf�M��y_��Ң�'/��+�m!zFgqY��f6�<�پ.lv`�O�I�:��u�;r6-��s�q����]=�Q��!o�\:!��&��aX� |��Z�.����G����:RNc֠oq�&Ѱ>��Kڶ�`�8�Y83�i�<�Nx-3�L���ɞI.��d�
�ط��ܧ�h��ߦٔ:�{�~o=ab��֐칋�9ܖZ��'�e�%VR_X=�o�@��<���?�K�j�nGG�@mv�#�����VN�.K啹�O�����Ŝ"Җ�}g��]x����ouj�~3��k)N��$h�:}��c�-$�X�_
�V�S�Ң�RZ�|��!Pzt��ކ�i�Xi/�01R2k��:��E�WT��S��.[�R ���x,U|9�R���|o��E�3,N%�$��m�����K�r�j�	� �\�˨5@��"�Ē��P��m�����=�Iƨ~��?l���#���˓��IN>�&yX|�i�L��٫�ܢ��,��2����<:.;��_�g�nْ��le$����CP����ko<&�G ��9��e=㝔��?x*�/�w�㓄5F�a(Y��3~D�>n`�i���g��L	���?4�9�}�8?Xj�/��+�`!a��l���c��:��u�D<nES�c�3dPKH��&��w���H�Y����3�
}���sO����>����;^�d���'�sS�#���� ��@K=*��]D�ܺ��R�I[�ys������ٱ�L 5�ޮ��([�<Vq���A�V���Z�ֹ���e���w�v��X��xeu�;N)t�#mb��nF����t��-�4%�4�Wϗsãg��E�t'4h%�1\(	o&|� ���-	���Kt�e��?�]ݰ��CEY�"V�I��Kɓ(�2�9�!�Թ�:}!3�9�wK�Y��|�^����V�� ����