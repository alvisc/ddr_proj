��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t�������.NT�ɯQ�_�EY�����]|�=�Ăt��@��{D;ӸBr���J��;��?�͠�j\i�ş%m&j��?v�W���tF��NO1���?!T�Tg�U-�(�	Z1��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HCZ�C�Ru�����[H��22P^��{������6�a�WN8�L�u�E�>F5��o{�R~�Y\m�Ȕ.��K�Q�ց2.����/8��cG��B�+�%Y栠��'ޭ�--j��7��ml.���~j�n����©�kh�ؐ��=?�^J.W�Ս�8�"n�B,�U��,�qQ�0��'vI�?�֐`6^�fv����x�Bڻ�.8��9X\�7������T���Z��َ
��2&7�g&���:�A��˝�9"�&"6("����6�4Q���ܗ�^Q�Πn�V4n�w�<|% ʨ#�p׾�=���$�&����p���̅Uh��/ʨ6�+�]_� <�E��3�?���굶�&�Qg�إ�ɉb���8k�a�\I�q��V�	�؟mJ;�K�&��X���n
dn4���^6�Ӎ8�%��j�|���uC��vQ�n�Y���5�B�|�:���zp�����cJ�[�}�|��ܻ�:� ��>���+ܙy�SB�+1�Fި�ۦnww��sTPo ��L��:a���V�:��.r'�7��⑬fY����{K�|"ra�өW�{�(4�kIW���k�7]���':��Y��--r���jɅj6Zi�LW�ڴt��<͡��i�&CX04�Z�S��H�R:�6�`�-�|*}(�����S�Q����W��(c��d�4�+32�(?���yJ����}X��7kp��9� �p?���Sޱp�gIq�Y�RҖ�hr3X��Xx6Y��p�Ϥe��A�� ))��L�nj���ǰHs>���ѧ�U��Ѱ�31��iI��%��R6*�^࿇���Rcg�#q�Sj��q�����s��+Mz�K0/}���B(@�Bʟ0�H�`h��qX)��*S�F��vn7���]�&g+zjѺl=�0�	���eW��
��tG<���m~H�/P����y�ءv�/ܙ��;�T V�|����!�F��#^���+k$��AR��qBg��e�*_�3=h<=n�ӂ�Y�@�ڟ���0�,{i�ybĮq��9�������L�dkL���[�S��B����v�N3�_�q���A��P9P\�.�/&>�{/1Ԁ�y�	:�31"�ϰR{�P��c��^��@��j�veJgH���3N4RGh��ƹv#)l�C*#A���ZK��#�C�$��Z��ji��Wy�T�B�@�4�2�Y�G����<'��J��@�&��|P���4�儌6Ypp��QBtS��B_j��� �y�8�o�I�\�7�p`QT��3�O��nd)�@��1&o��0rbT�4m�GQC�����\�>��|+|.�n�kI^Z�ǿ��ݕY��-[ě�Uc�k�! [�)"�ٟ=�c��<<b3���� ���gv��h)��*���V_C�_GA�oѽͱ-,�)>
��q��xvt��˧�]��-M/ϧ�m§УlF�E b ��6Υzy�F-6�Y$s
�����Y�x�^$q�ew�U�r��8��O�������K(.��O�c�}���U,��Tʃֳ�]�B�nv�]Ht�&������@x��޻�W��&��� H:5���c����k\���Y��N��$B�%�!HL�M��z�g���h��k<oM����вjNGl��f�#����Ir׶�1�q<�	r�Ѻ
�<�a�^.װ}��)�h�/X�9�$��i�\�K�ަ
�Ւ���M�F���<b"�wE
	�'�����q�hV5xl��~��'#4��Q�L�0'O�k5��J59�Y�R��6�������U��x,�7Ws��0���s�a�x�Ai<��璹��������C��W���q�^2S���*�B�0��e��^ӯ��f7��]� ��m���po�~iG��4L2�?�y��zW�+�:����I�
�ct�y�%8g� %@Y��rx�*7��A�x�7T���6K�u�#�N{t��"���~6mg��3Tw/Ad�_𫳑�����%��E�4^�Q�U�7`Mx~~�i�һ�=���d2:$�b�H�IB�+��"�0q��o@�x�_�o��Nr�l>�b���P�!� 	K"0'��C��I|�@�v���|uJ�,��07.��7�n[�1�քR.!����o�.9;9Kn��`���@�Q:	К�#9�>��34M�SuX�c�MrL�W��ځ{����"��=߯�Ԍ��F�� �DM
�t}r������t[/��c49�c���c�h�N$0���{���X�fg]2��`X���#N���=][E�܃R�I�z��o!	Rtկ��cѭ�i[(��n��B���	s�9í��T_�ܥD�>��Ʊ�Zp�^[R
��1!6�{e���,��|�;�,KW��lڹ��)���`]�)s`��!/�y�ޠRǟ�^s�S��Zʜ'�<���_����n^Ӛt*�	(ٖ��	�O�����E��z�H@Sp�k���r-�~-_l�`"ޖ���u�{�h�;&��Tp�g�vppƿ&��a�������!?Ա�N�6?iT�.�ja?�G��~������`: ��'�=]��T��������#��4{�1��im���� (���y����O&���Ev����J`�8H.��%�K3DM��&$^b�I�'xݓ(�X��9)i+J�i��8�#�^��*�<���ˆ��E2�z�cԅ�O̞5wj�� FŹ��O���Kg�`��_�NҢ#*�����q2{�$\{]���Ś^l|�����!?�8_y����@yj�RϾ><�>��<���m����h,�ey}�\|���������\W|����(x8�δ��\���Q�Nz��*3�BYoTLp{�NsUo+��'��UG�Цl[q�Ƙo�	���~�6oFٖ��a�ge�~�4�tCw�2���I!�XX�e�A䤝� �O�u��1�����eUzJ��nB!u?���2�H)\~d&ć;5+;�㱧�"(A����}HWݸ��M� ���ϱ���uHт{ȥ�"9XV{5Vs� i9>%,��O�5;�7�Ǻ�Hn�<a}T�ߥ�S�|�􏡚�G�8Z��?3q�ī�\0r`��gVE�.�yFyhVK�q��\��������Tl5��֙U�nV��X�)Y,~���'�F�U�Iױe��h��u��l�7���MF��P�A��Mkn�x+��*ԶsPB�bg�&��N|�#��uaa���M9���k�����;�4��l�iT��Ӊ���I��XfvKO1�3��[tN?�᧒���H�*,G�}�<�;PaDF��J?���}I�Sח����0�Lt\	����y��BO��҆�|��ho�H�����Jp�S��М��8c��|���h�n�FC��.�nv����͘��N�l��J�S��P�ϽC�IP�M�n}֊�ѻ��XJwK�Q?�Ǆ4� _��2[@E(Ŵ�=F��7.�Xs�#���%�q|��y�b�NV%���Qǟ3��i�sⱬr�	xͽ� fi�9I:L��ԺT���%�ѯA	�-��}��R�Q�.pI�B�?w�K�{�U�b�ү=к����]�m�H�}�E�<�ڨP߆�X�m���Va���c�&��O��Gp:�36o[��5�{.Ѝ�B�~�&��LBe��x�ǆxsi0t"��A��� ͏��63�k�J�y�Qs.���<M)�XT?ܦ��<�G��-��Т��k�����Sƚ���ᴤ��ö�9�� ������[�
�ː*]��Ǥo���B �~��`\(
�rYuTN��}�8N�L��5W�%�Mi��]!m�*]���l�L�O��=+�Ѡ~��t���n��Vg7-'�z����@��P)e�ݛQ1�����{#3�.��k��兼z	��C9��pi�d��� ��ьl�=]b�
J�g<��l�7;�'��E8���-Z?�h�	��!��LEIF�x����OA�i��S7��f8��>m���+֔q��Z��T �A�F��Ы�V�'�|À�h|]�/�u�)���s��~���Clf�o��e�mA���3��������m�^��l����PЪ����������5Cv�t~��k�q_5�4�#�	����z�|�*�ѡ��]��0n��ɶ:3ǭ���Fα�Gd�o�0��=-���E֐A~�{��ސ�� /#g(�*S��S�O�3=�/#��C��2�Q{�<�Ӫk�}I"TNU�Iw�$p��(�a#��*bs��*
m�� !j���M��H��a� 	�4Ӊ}�^�^=�!w�s�-U�Qv��܉�)�q�˵/�W�h%�1��6Fvr�S��ֽ�F޸�9 �`:����#d:��Pŀ
��>Si2ǭr"�!�f��[���l�
���0�c]��/)�<Y�%幮����3�G<�R!6L|^��VY��o�,������H�r�{�g������O�F~ؿ�7 8] D^�qe��&2��|�`�񥫶f�g@]�YY���^	g$<JE�t���O�ݒ�I�s���L�?���u���C�=I���Sq�Y-�R���t�v�#���B'"R�V��!&�����m�  W�t$7w����u�>�ϷR�6��������t�_�x[�����;������t�6@��&�a�K�K���ۯ?�1�|�r1i̐��S�f4�F�o��������]�~C�n$IIµx���&:r����&a��9Ȓ�����Tj�?B
Z��B�\��ȫ̭��ߘ��F\j�q6�h�4��bI�v0�&R,�T��ks��}7��ўa[˧��ڈY�عтb;���
 ����d���4����O�[���:�'lB�*�v����j���x;���p�"���)/X<��U9Ԗ������=�O~�@�{�n�S�ǖ�􈱮�_p�v��S�3ej4�5�Yk�
���"��=N���AI�i(���Z�-\J�N�N&�mcɀiL;N��%�,QB:e����:���U�I^�l����=�#^��tM�8Jᰍ�O��p�fj���TU\z
$�m��ܨ�f����Bs�|��|<
����g/����9G->�q-BND�x4�+�z���;��M���
����&N%6���P2�S����>���IJC�v'�zk]^[qe��\���+�DM8�yRޟ�l��YF��۾�?��$��)B������D��P�}�V�\<��g����$O��Ң�>�v�b��F�οG���B��g��|�hQu������w!�e}�	M�63/2�.֏pL�d_��]�X��d�������<P�����A9�7��љᣈ��*.���6���_�����c���$���?�r1�d�	l�9�Ƙ�B����RVv��8���V�0��jsv#�ט�L,>|)�"4�>^��v{3�5`P�+�a.��,����m4������A�}'$H���q0tY������|ۃO���$�IQ���z%��n6��3�Č���a���l�ad�|���s�~�6l��@�GZ���.�g��/�7���p"�BU�hH�Z�֎z��������Q �R��Hu�9u����m�I�.X��(��d'�T��+���,��Q�h��B�S�v����#���u:H�˙�/��H/�p<�h�g��/�("�Ly��ӏ��?�/���4�ă"�2&�GLSŰg"BZ��w�`�,�� �J1Q�]�)O]�(�BOf��c�R�xq�\s5���)�\�<��q�"��� ���F�@�6]���(�;N�+�\��ξ�%Zg	Q�P���UFH��F	�n�fm���1.�^�o�s�:!G����KF���ʓ�j��W�z�F��X���(��r��ᦑ�u��K����k�46<ޜ>!�s��n�ɍ�4�M���<1ˤ���Y^��A���̡����A?}�qx+f���Ԓ�]�����+Zi�A-Mr�p@�)�)%��s�v�"9a�+'�['�� KK7?"V�����"-W��) �-*��T��74�k\t"xt�	t\�O/%�NLaXwnXf��bY��5��? wW�fm�n�%���Ի�S�4�er.zv�\l�v)8@˧�:� H�Q�L��������p|�V���lA�eՉ�pB�������A��#1fL�S=b	!m���U����ke�怕��}��>��X:@
�$�*b��)��K$�eU��2༾i�M�v�hl�p{x���e���-T�qY#I����h��ɞ�;�t�a3	Yťƞ�2U7E��A+�k��<7�TER�ͺ�#Xi�䙐^
p���vgF\,�,B�Kԫ*7��2�e��-o�*��`$�Z3�%�����
�b1FB��s��k�u�"kS��6��S/�{2�F ���6�
 E�)Eo�z�.־�����DQ�;Hx;O�"��*5�v�	��M�]�r��b��X�~�9t�ʁ�H���o�ò�����V�s.y��4��	uǬh"�w���0�)�%˪x�@\�U]�s��*��H2n_"1C��+���:��W%{�*L�N�P����� �,�ǝ1��Cw���v�E���j�oh��$S��f�D&~�
DHK���0�ǽ�[��1�6��cP4��/�7F��B^�����,�D>>��mӨV�_��E#��Z]���̰!F�Si{�F����&B�U�Ա�I�D4��z�	Q�0��������,�5�w����w���_d�#�v�]?�4򀻽p�w��_9á��A�وĚ(��4�h�O��G�F��W�8m] ��Ofυ�f�>��V�L{�L��8��UE;D�y��{���i�ؕ��)h
y[�U�ۖ4����x�1F�}�n:h�ҵ&�1�-���ެ� =Ә"�z�V"��#&Bq���$(��y�(��0����o�
�)��!m����a	M�[xa��i�,�JWlYBW#�W��+gB]�,X�M�&��R�=l8V�m1�h�x�=�5�x���蘦yZ�:�)����@8��}I�u�2�5���??����$ǲt	�\�	�'��\냔�XL�b���480�G,�kl�C�w�6z�f�m�^�S�	�N+0n4q�p��r�%���.�B��E!��4]�s�P_�O�!z{�4�7�]c������$� @��u;GB&����S58�S��>���WR�@���YX%�Xx��MN� y϶y�Ձ{�u)k��>h|��c^-�k]^nnrEP YZH�=���Y��A;�֢�(^=�-�2�B(�P��&+ed�����|WzƦ?��z��>\��x7
m�RyV��_p��!Hc�[�v[�
���6''�~�ѹ�H=\]��#W��F5�x�_6�e��zHyJi
^�a��ì�V	�edEƽ��n�n���3��b	I�F�Wn�J߈��dizu��;+�ܲ~l��V��ڨ�!�a��Q��w��}*;Oƻ���0���L�B������� *{l�M�,��%B�4ݼ�Φ=T�)
(��`��KiI�Q2������7<M��v�y8�5�\qP�u[T%$.=*ݷ$�G�|��]�X�otIca3L��?�ٴ��K2E��rO����m,�S�kr��WXB�`�s���{Vl��cs<Z�V���K�VG�W�|�In��.T�������s��A�����XV4{���߇���dC��@�oxֹp�e����opSɚ������o���Eݫ�}vi��GW�J��n�q��#������>w ��[��)�R�!5�3�i>g��O������'n��DI��٢�L��6���� ��e�˽γvtՉ�H:}�����O̧��W@c�g���S���t�L'y�b���\�yK��=����2iΛ�y��D��׆�;x=^8C��`��~w���lW�����u}Ss����F�#����\�X��*l<��)'R����:?H��9^�\�i�k&�U%�ఉ]�~G�k���ZM��S�/�Θ�΁qse����Z��!�����>X�*��OŹ��r��o�X%�2�	���U>���}�����&����ڋ� #������k??�
�@G�.�Tԉ��ד�����M�ǐ�Y�Fu�t��[��9��Q�sȢ�B{ŔNl�dd��Iϒ��[)B���ɹx��kd8��_m�
}�*V#ZO���t��$��R�a��� ��Uxf�r�q��#q�2&!�`l#�aDɿ9��������}���>ի��L�������E��K]}�%��B[�v�
��c� �Bg:�w��r��^c`��~�U\�@��P��v7�q��X�nyב^�9L��rg֜�j�d�^�3S���1�y��}�ݱ���YO�A5+N��s�����$HR���V8K�Io�E��D
[�-Қ�$�魹�=-:%�*=�P�"���ŋ$�:�|�a[�r�v��-�1*LU��7��8�)�y�,8�1�#��M������Y\��q��k�$>��q`;�gw���7u�)p�9��#޲�c�rbRHZI0�+������K�l�#��F�)�^&[���
��wI�sxK�to�4*r[���N����蒵�W*k��Ђ��}2m����@�h$349����c�����/jJ�z(C^��W?{Yfx���X	�Y!'q�B�N>��Xӓm��d��o�f��J�t<�GX����R��>v��;iR0����}vdV��`�k�!>�G���0{���61�T~��)$�!&�����{���)��qQ�-yٕ�a�@�w�QH���R*�;��4��ǲG��@:l��mq�E�P-9\�*w�����&~���{�G��y����V��D�݉y~휑����_���SK�0��.2��WJ��ǋ/���xz�4X6XQ���,aB!/
|
�2��%h^��d���4|8�V��b)=�����>C7�D�O?�v�Z��fwV��wї���%�]V�^�	��S�>��b��[xC���ue۱�M��>����ůuM!*���Ւ�H�����q�M!��B���N��ج+�����&���Ʒ���ڸ6�� ����#�5�UN��~��t�Z��N�5��n��z�U��vZx�G�9{P ��N^�p^"�/�Z�=L\zB�o��!r	��]�ʌB�A`��31C���J��~�ȴ~�d��~qT��wR/�"����ڊ|v9*|љ�h*%�����6�U��%��O}^�n��J����?.�&���J��ɛ+���R���ѷ5��}h�#��'�h�<��N�[�F*�q0i�z��C�1�/�\8���f�!_��6�>����>�*)� %/֮B -�����B\ �|ş�B$Хư?�`����) ��o�H)8a�7O_2v����q�M��_6���;�)Qk�s�����i�6q~�����Nn���	j��H}�Y��Ƹ�.����m����}�w���3��`���G���}�ȝ�kȕ<D�A�)(�J;�Z���Rj�1�<hZ1̒",h0�o�x,�ӻ#�vY���1(QI^i=��+�~���4�ݿR�|y7}�X�2$dz���p�i�=c�f-+�����y��Kn�o�?K)&y�O��<+cQ�nЩ�Ă�ȳ�!�;�����\5'z0�y-ˎ)�蟧!��]�_��X�G�ih��E�ӫ�Q��M��r���+R����(�����n͵�q	a�%�Vl���:�b� �2�&?�1G
���c���٢I������`}�S�P�ya�G9��(� +	Q��'-��^��l?������~J|��~��&��Db�R��|��tu�����U��l�lx��Y�>.�~�g��K�!�(�]+MF'���<8�$��h���Q�$�n|�cv���~m8=:��\��3E����ۀ�.���NsZ�c�\^�� ^�{������_˸{rn|�JQ҃O��P���}�|n����-Nm��5y�e���c�Db �?/���Y����(k�g�����;/jדo0�@a724����е>�a_|&
ON۾	�j�j�$v?6ڃG����2�n ��ֿ򟹒U��Q�w^����v�I� �RW���������l�~��_ V�}�ۣ@Ϳ��w����������JK������_�U��Y[�8Ci6���|�Ppm4�[�eX1Gb���dq��yMXm>-�kc��~v�*p�X�ݩ��2ea�Ã6��6��W!��6��(ā�cu�E�f鸎%����Yn���M/�F1�ӡ,��-*'y��&����*�&F]�K�����z7�(���N����:�v�@�Q��x�i�C�|$�݌2R��3Q����\-(���=�J3?���gѺ�%�T���)k�U��s�b��0���Qb����_���s�)>�����#N�����)#�]�׮E�0x�Ύ5�[uj���i9~�����5��b�����v���`��ny�t���*<�ɕ}$sն_-������k�ŏ���ȸ��I⒤���c�4��m���j������~��:ΝI�˪�@?���3�!5;:�)�� ���il,�Q9�C��&�EhA;�V�^f��׸�E�ϯ�eR��W$ ��3�^:��^�L$�J��$�`�_��� ����O�bHbX�Y��"�@�=�!��i���{����5�v�a*��Bv���=쇁Z%��x�`��p�U��A]�'���ZQ��is������q�%(�ާA?�N�z���LF?pP�Y���k��d��qfB���9�z�zH�:?&64�;Nxx��O`_=dѾ����z~VZχ��:��ü:F���^h�nu�Ƞ3A�12Ys�6<d�,QoI~���[�]5�������|ir���2��ܺ�&�TL��Ͼ-��d���<��[�:̲������^�򙇱�N���dR	F8��C}&yN0��������<��~Ř������nlaP���kg�����иv���R<�+`�e�H��a�'��<��3G].��j�p��-���z\�}e���q�򯡎���h!�ɺ^�Km)4B��������Cq|)(��;J�	����p];���1�9�x���Pi�$���Z���W_0Ť�k����+?���<���7���^_����!Is9��3���1*D�;Y�VU�ֱ�}OQ����#�N��H�o�'��������=�	�:׿=	I��1�	�G��$EZ�ń�{"�?Va�%F����Y��u��[�,{>I�BzV�\d�9����}4M\��V��9�-��-!9�*��Wt�5O�:�D��6X�e�O�`Hue,��&���9o�ֈ�{2���FM�#M-�R9Qr6_�I���e�Lw�%m�jhɺ�	q��\*���*�A��̢����z����	����g��< tY竅r}@�Vv�sd.��u�	6ۑ�gb�:ԾAK.1'��I���.8KB��ݏN��:J(-��du��5�����e��:%�fT��A�g�!�)L�W�u��5���V�Q{������3�!Z b�~�lo[�Agyr$5����QB�>\��5�<q�E��/~��O����zm�^�׷���ϑ뺣I��cf޳i}���H���{OR�m�Z/e�!�.IgD�N�ɳ�rk*�� q[��K��bk�N/�X��K(�i�6p=�N��,�I��M���n�s��b�JL����^����Fd+F��[��u�o�V͂bϊ��<:����0�>���g��f�@��)4�KOy��;��S2����KSK�hb/���\\� �� Ȫ��
D�K����j�`��Ej�uM�R���_����	�"�C�J�
�6�X]��[�-��z�mߟ<!�!�Pa��1�4q��X�mۑB9�J����f�r�608+�c5�k5x>x�R��¾W�����p����쇩�޽O��O>u��UGf[�Br �RאZ(��^/��	Ę���5�@��vuuH#���N�5���j��-�������z��!���-����L�����/���c�����hm\���~g.x����#%G�g�����<e���H��N����/��[q���j���V�w����/@�l;��-��\���[03��o2i�/��1_���B��7�H޽�����ӾS���1x��W�)"~(h~�g�x��,Id�p��u�0F�L>�K�z�];4C��9f(�&��C�2]��6�q$ɍ�WL#��!��!af"^�U"SD����ѦJ��"\V�'�8t�[�rC܀��8�r�$6��!
���z�X�����lO�3_�������������ဎ5�`��"���M�S�#_ ٗ�HGBh%A&'M�T�}�}���r4�Q�]x~;���5q����%�S�%��8�`�Kbi�y�H���7�P�e���8������`Q"�ե�{�46�S��a)�36B�_vH����@5�O�44���=�$�?bݴ���
K@�kj�U�;�fǾΥ�Sۯ�Q�&�A�α��,R<�H�v���������&*)hFri�&�͝I#ϋ�
�Z�����Gs9�J��E���I�ovpSd(X&�ڰ=~��o1ޚM��CD��~j|��qA^Y �>��e��<�t��WI�I$����E
�
t��O�(��A��6g�i�*��_gT�b�mZ.���g��Ϣom�	���%3DG�KX���VF'C-�a/��Z6?&�7��Up�@{~�7�Rݖ�y�������b��F[�C�
�b?�ģS/]�Nk�� ��Zۡ�β���+��"�r����HI�M�yz�ߣ��R�́����'���I�{�>Ҁ�G�)�͗6�\��Me$w��M2�����J#)�ĝ�ȈIz�]�c���9��L
�� Yvƞ�%���l�F�i�$��^�[3���?k���#u�Ն���Iɰ�^d{��h_���������\��R�l�����<ZK����ƕB���t�:N�V[�s�}p	;mKжȫ'|%ӄF��2>F��܎���\X��w����5a�3���m�Z��ٔb ��=.%���9���?�w��RK��4�P'l̟�龷�]S��U�ݒ����=D�	��nCa[)�#0e�+	�F6 ���d���T��8���Y���M8��#�
��/�Q�:�B,��&�YK�|*5ŊB�8 �����P7'�a_���*�>W�`����+F�go����u�ۺ���CD0{ĒSڝ�%����s�$-�<>�NtJ���J��N�hN���#yN��4#Jf�p�D��-��/���(?�i/���? �:���t,8u7%,u<Dxp1l0��?�YBZ�xc���]����Pf���V�<��r.2p)��k��ɰT�{gS�8�>�=Twi?YH������PEQ�0�p��ǧ4�i�]"��vGw��#�#}�rR��\x:�M� Z�?z�N�A��U%����i���|�^�VD��D��~��S�b?-�����j<����f�ܩ �8{��3��|�]�?.>X5=&��&%^�\���g ��Ȳ�+}��⚶z�G�	T*��	���e�Xr�|��1����~B�gv��tq)Q����s�auȞ��_�b5-٬.�|�B���e�� �d1�P��aj)�;4�[�U.W%#'�1�<�{V$'�w�����^�vtX-��¾���Ū��9�}"���_�'iI;7��D�EUNɈ��no/ȼ�e6rц��u�tb"�$��������H�p�Qg:h��>���8;�@�_�> ���� �`I5r�ۘi��v�F���
��O�`Z�a��*�������r��:G�p�A&L��ɰ蘙%t��N�1Go��)y'&��β�w���b�2w�Q!�x)W�A�:���٧=\e ��c�@�<�@}C8��#}`Sd�I���"A �#5L�lG���ѱs���|X`We갓�1������ �Frs��*��!��= {�T���JCH�R����>�����>�w|�%7�^4bM����(�XBL�G��/]���E��m��6����
6�	ɦO��Yv�T7:�/�7�	�UAU�"%K�����_�5壊���e��Ox(��L)6���p�K�H�nX쨭Ua&RםG-�/��'2d!���vE����]!L���`�#`h+�q��c_@�=�����#�\EM��<Z��> �L$��Y�i[�e������\���L9�]A�0 �f�0ʻ�n��w �.�������H�j5���MJ�!j�~���F�]�)�*0���)� �,�ui�A
M�w�em����9�j]7�7?-�_m
oZ���=�K����)�5���x���
�i�"����R�=n�5�  �T!Wb��/���}.<V���=ҍ9(Ŗ-���~i�,��'�*T�p�%;g�8J��C����l�\rM55�d�9��A'����T36g��9�񕚍g@��q�;l�8l�Fzo ^q�s,�����}�pny�&�B�)e΀V<�J���	F���X�A
�)�<K^h0hLϬ�VB��Ѯ+���_R����l��?Z��z�L�|���T��.�)'���Ă#�X�!7��rUe]��9�n}�Y.�Pn�����W��EQo��|�1b?׎~��A��=�_��8�w�+�H��
:��Y��!��=��e3']��*%6��;���Q�gk�<��G�����!{
	8�c��ˡ�G�h�Yƭv�t� N�RF�%�|�))��_Um�;����r¦��_1S�_��絽^��X���%Y�"V*s�3�Lw�K��44�t��~[n����hɴ�6%ܭ�(ӓ��.�I;
����SY�k#$�ś�?���Xп��za��3��.˗̵����Ț敭��d����jS��q��\@6��ra2���˾�x`Kz6�ə��m��L�Ǚ�jW���@M��YRn��>l�3�i�׸I�'vc��U�a�s�	�FS��f3���=�V_1�TF��	N:��ִ��[���L��`i��Ma�g�� "�'ͽ�4�h���j��f�r`��}�������J,F��V�g��/�E��W�X9�c�H�a�!-
�;��Y��pQ���K>�s�h]3jG0�(S���xҷ~��ʡ�>�"�Ee��lZ�kq�V7,C��tnD��i۰g
Lk=���k#������uR�-w�;�-v����gC��U�,�$ՠ6��P�0ڨ��k��n<���f��H�zQ�`�Դ��q�������Χn���?*����Z�"C��$V��I���Wg��q�'Y����"�lbp��{Y��U�P(�*���K�r�%|�Snv�V/�ÖuW���7�=�Q�6��#(8C����80��
�I��@��n�I#i �[�`j�2tr�᭓�-�KOs��zf��ݶK��IS��es��g}�0���K�����!M��W�Jq�AA�P�("ɎH�G0��w�t��a �+���;��o�;�Z��em��"	��z	��n�V!� �U^��S�����]E@�����&)��2��%l��c뼜��@\�=NJ��h�8��Js����[+t�����+�+���]��*�$F�����`t�w�)�$ �w�?GF��o{:m�b6�Y[&��b�	e�4�k\	��LҨ��!�O�Fm�Z;��ƳIG�I��AG1����/5�4f5�����]Tmi��(P�z�Orp�zME')ZCy׀��9�µ4#��k��\y<��o �[�KT䴃��F��+�GE��H�5��X?��G� '��%�Εbi�e�m��n�rq�,
R��n%B,�<1s��l5��
uN=;fG^o'�Ҙx�?V�QO>��y�3t�� �����]�,@�(	�Y�5v(��N���Ǆ:�F�4t?+Ӓ��|��{�cFh#�RV��Y��zT��e�Į�|��T���s����4�{��B��Rr�o��㞷�OL6 ��y�q�Z�Waj~*CE��̊(R=[]�L
:��v&�k�v��l�S�MB�vl��W�d��p�"EmU�����KARYc���wŗ$|�`�deF��LƠWk�&M�̛N�8�<|�T/!�F�?o�{�}7�mpjqz,}
����!�f�w#�PG���KJ����U�`ȷ�@".�]��k<p��S��U��Ɇ�˽#�ی�+E������^�Č�r8��D7q� �Q�Y�����hqh���ݐ�%�@VH�6������t�r�Fn�U3P�?h?�c�����Qw�*-����Ӧ�v$!���D�-�P1�!�2�ɿE^ p�/L�����O�������Z�vhZ��ŨX�D�{X�Kh�:
��z�Ae��]�g��V��<���Y7}��K�SI$� _�
���m�&6�ҋ|�����R�a�������R\���+v��8�ĪT��	�PF�8��+�з���t븖���&|��,&߄C�ܤQc&���I�gY r咪�����Yh��ho���^��v�zz߇P�DB��:a+ì�f!��P5�tl<�K�P�Н��I!М��i9����n��rQo�(U���)�>Rf�(��?��!*�^��Wa%z9k��|�	X�ٰ_K���E����p��9�A�cm��}�Zm���"��Sm/�?��f�R�Ҟ] �;�Xm
qYs����4 ,� ���֊��q��٘��l�7�eS��r�EO1�p��f�uߕ2���*�@�?�p���Xt�Ԯ�G�ڤ���?�Xf����,�"�CC���ը�a�T8�/���5�*��,��L�SV����b�}oZ��c'�GxT��� ��l�Y�+�a�uގǲ(b}�c�Q�!��ʅ��c[5SOC^&$&iv���H�8RU���^Fq�3�Sn�ϴ��ũ�p�ҡ�uA�J]E��C���=�J��a'v��@r\a�7Ʋ
<j�Gt݇?�@?�'e��T�@l�Ѯՠb��܏��R>�B���ٜ���m\����1��/�# 
�m.s��~�r�Bb6�i;�F��M�X���F���KT�%
�s���ϐ��MnzL:����<��4��<�͓�O^���B�����G<�:�ɠ�M��ed8�:�V���d��#Fp�Q��"=�4UI�zFx����J:��,U)�s _�
F(��@����CT�v2�R�
 �>X�	���zH@m���p�T�S�a��FJ�W��%�)6�z�����`��{l� ���i�)����R6se���Ʈ����XB~��1D���;pkE b!���J�=X����gVќjع����6��!���8g��?!µgA��H �����1�7-���*(��d��cTS�.��V����C���� }�r-M�{�s�n�3��0��[#��dD��s)�s��C��WA���>f��Ӌ��C+D�%L���ѝ��K=[�J��%�[���m��fִ6^��"fë7Y%se�7��
'�R�hEO+QD~N�F�(z��v�k��s�5�}�+�M�?�� wɢ��O!���	{��&l��Gl�_����z��P���ܘ�����"�v����m��Z&$�k%�K�al�J���$���Ɖf>D����IpK�]�x
������pڱ�TGV�r��$���[���R����)��<dK�C�^�}�l�V]�y���8寯����ëa8�����؁�P�0��WN6�B\��<����Y���j��Q�o��ũ�{JG;D?��6ti^��GYg�d��_�k̂��O�d���7I���]�.>��z��V���ᇿ݋r�a�?8��iNZ��=�G�J:�U>�7ؼ���q/8u�jУ��z�h�jv�� ����QC:09�}!�[-���S�����Yw�_�2?��PV��-#�<]ӏ>�k��s��)Xq���d�C�*�v?�zg����@��/]�sN����l�~��"�R0��/`s��56Ty�N/����ݿ�҅ڂ?.F	�����'�	R��Qc��^�g�cڍш�礆�Ĝ���V,��u$�J�|3�����MB���/u���Y��p$�i�
�3��2�uP2h� � �,9G/O|��J��7:�h�n�8��ɷy�t��#�/Z��k���qS`;?1������H%�cZ�)h�|�3�ȇ�b�p$j����W�<���g�.N5���(�m�Ѩ�>`e.�3����b�hD3�s�;��r(����^3Շ����SN�Q.,|����Rw�M1�� �?3��-�B��5�+�����r'KtM��d%��30Զf��m�.N�@Y�0����[?��X򬿵>}F/��L�*�.�E�ȁQ6M8Ru�̪&��p���6�K��^���	$q0ie/-+�_֦�O��n�)�.Ţ6
�ԏVG&L��%1͌�5�j�9�9����rL�D��Da`T�i�8�?��I.3]W9�]3�^�A��ke>�ONșU��$��E͍ 5���f���J�"{���P��," A�2��B`aC�j!����f �����.u!1��7c��y�(W���ra�L�w@";�n���o�M�
�].�W���`�8�I���Qr��i�Џ��p��5��0v���2����v���+��+�Þ���O��Ő���H�ϴÛ��+{e��R�l`�T�J;m7�)	E�nAfM��������W��{�wpZK�@H��]�
�q���,-Kp*l�^���jc��L &�w��ڿ��iu��@@��y�����>VPE�생<���  	��	C��au�U(�EEV)oh�>(�Ax�m	��31X<������b�teIP�M*"w#��i�g�1�eҪ �[�:5y���O�k��(X�Z>����Y��E֡n�bLM4�"e����J������彥��b�B�奺�Ǫ?Ӵ�q��h�/���f@�/�]GF[ ���M`���[���Iae̷�v��7d~%y���y�B��AˀS+�?�ȷ��XJQ���il^��lK���[U��&̘�5�,��ɿhjYu �����j*0�����*�b5�:�����ʛj��W��7&��E�K=�.W8�4B�5>I�g�"�_s��Y�����X���:�k&�K̳L�@��5������� wJ�0�U��Rw����)����ql�l�b�S���������و�#���;�I|뒊yŦ����Ǐ*tڱ�&	w�3����.��C4��\
����nP[��_�KQM��oI�cHM*�1}�!�!�j�Dw�,�Uj��BX�E�?Pg;d�ms���z���\��q�����nG[�eLl���c��������L�5�[} ��Z'p�j���C�,a/��,�@��>�" �tb�'����dȻT1B�]>N{�d�����ҥ͆���ĺ��E���{����pp��Xl��B�D�|� m�9�b	�#>u�C�Yf�'��;5�^��Rp��k���<�}>���n�ԹH�Y�|&?f|=?�<���me2��M9]�b(B��s���> )���] ����?;�h)�5�8GS$�:Auܖ?{��;��k[����L������@  ����-�LB�p1��ͪ���zxk�3/�bX�y����^I��ݠ��X��ܧ�P�N�H��!�\�D�^r�p���_AZm�?�����d ��o�S�K<�HdP|M�X�+��A�kO��|��CȞ� sOl�]���;�Q|�:��`��"�� ��l�K�������#l��a�0��0�R��	f�Z,di){��uҩ%�zP|`<�#:�B��u�S�3Y�bQ���q���^#8�������4[������Y�HO���@��/��З__��+���(�7�R��*	�fߌ��_�(}��m�A�ܑ�GΪ�J.�>G�����q�;�<��w]F�r�ط�@�:Z���N��=~���5��"�gzm�0`�C3$~Z�:E�����f58�����%K d<}$i*�š����YzH�A��xn�
 ����U�˻]&��џ��
��
Mݻ�H��5(a��]����i6�jB�$43Y�F��Em��_�ǯ���ja��_�Y\����8๓�o�G����U�{����ݻ�~޲̉��q�7��5m!2�׎�,���^�Z��:k�)c�e^���t�
����({,���:�bj�� 4���7�����^m����\��x�]Er�]Jۉ~�׸��81�]T�V��&�=�u�\� �v���sC^�4[D�Y���sk�bmm2r��������f�˷�?��f�2//��c��e��_�ś�v�}2�R�|;�Qr�}[Np�}ҋ�����gJE�m�e�6t1�����d�G� �e�j�4-�y�3���_0n�~7 �޼�����v����}Rϟ*�c�<z�e��c�So���w����|���l�z0�e�g��'�����	@4_<�HS�OV��$��z6��o�J�*uq�Z�f�bM�F#O�.��N�j��'��N�⇑�5���́-��aq��o�� ��n�Jh2��-xa����;�`�D��|�@����V�����E��% �7
�|f-��cTb��5�D�.��]X@83��R�	 s�z
 t�J%C�m�%���;��u�H�ݗ�� DC�Rf�#�*���,rfVq�.W�F��Ex���`&B9/ӱ�TE����Zt�R�iDJLO�lJ�\��,4��v���_Z����I�å��r�� �\*^�df}����!v�piߓĝ�����+i���@�~��0���E�W�yg=+E8ٗw�NW���␹�9��t�K����\�b�~
�2�)AGs���@0E�#3�����}++�9�A�dV�D�=OA�G��$-��?�	/�h6@5�4J0V�H3p~j�J[�߭h�&i�����H��1%�5:6jC�"��5>�<i�.D���'� ҉W0���w/{�*~���l��yP����'=+�W��j���^��`Sg�Pg��\���	|���Ԙ� +
F��ţ@��ro�`�Er�dw��W�
���/{O�
�����;.ͼ�"UqNs�+���,(
��'�~�[d�!�SeZ� �%AuK��?	2t��}i��d�Qn��O#�ũ	�?`�`�q%�[�T��g .��^lݬP�C��P��x3~����t�&="vR'p���:�"\(��8��2�A��6u�)^O��M'�A7����oa9�6F5D_��M^�irI���Gp?�z���;-��^,0��ނ#E�rj��R��w��������������9���L���mҦ}㚝7���d����%�a�J��ia�	�HoJH9���Ѿ�am�Nky��c{�����̬C,_ޱc��p&7��Ղ��	����@~}"L���(���(q��sO�^d����`���~՜���/m���F�U�_�H@���9RW�b~�-Kѱ�by�l`Ζ:����������r����|ʤ�SCk�g}��<l�!˽����7$��a砻��,ɜ�c�@��>�~�	٭�T�u62��cu�n�tO������Ҩ���>���"�f��/Q)g���j�b��X��R��Kc�mI ����m��{��=���y���߭��Qo�ˁ�6ǻ�4����\��,:�KZlD �ז��|@��/�AF��_j��0l�@�Hyu�7z~Xg.7H;?�18r��$¼D��E�Ho��a9v`w��!�	D������������Y�J�ῃ�ɍ lZ RGC��5TD'��w2tv����:~j�5�"� �M˽�؄���;�� Gf$�"�!��-�-������89"���4�92�ḱg�*PA�������9^|�ꀩd��Y��O�G��0>�B}������GDF�A��#�K�(,���,�{�-v_2e
�*� 3g�*O�&��o�
�q4�E��d�[:�3�V����/�M���LC��$�H�5Jy 6�C��e 64������c�gX�.���C6��e���MO$��
�jk0�-�5ؓ�ob���r��$C�|!W��J�������Oh���6mrSï	7j��-F��-1�(�t�G��ے��9��-���J�l������vX��<H��y�}�� "��2��?������u$��"�W{ױ�ʷt߼���)�v2����2�ŕ�f�TK��Z}[���a����%��f��-�k���%��	L���0�R&+��І?�^(��8�,4�ʇ��4��>�=��Iikv�*�ع?.Pg\���+K���0f�L�3-��<N"�P�q�|X��pS��_&K�FA������4m�J�J��,�M�yX0����,1��P�%$#�̞ O�3:꾼�֩d�N5�oI����1=�Glbv5�5���?ٗl��7᥼�a�͇��X)4��o_�kqIK#3�1�����r��x�Ih�B����"<\�uLAX��$B��n���E�\t�������l����l3$�H��*��r��k(ߔ��5��NE��K��Þ��	:�YS7��D�ɡ�0��1�6=j��)�cМ� �O�U2��wp:Ue�~���kW�:��f�%A\��Bb����)��4����#&c2��b,�5�����"�6��P�I�Y�5h��ީ��řF[l�Z\KX�&T��k�
��\�fkCD�^<�]�g�P��
j{A������Md�c�?x���U!�����V�Ym� ����_0g����k��!s�Q]��a�&;�I>eO��A����x�����Si,�Q��N5�����&2��>��m�!�r�tE��~3:g!�F�Ix�>���;���sӗ�6�5�.� stEC%d�lH�d��N�f&7�j�����d�T��7�W4��b��K�I�~��a����W���K�ՠL8�H���b��	�$bcGKP�&����7�O����4��|d���X�Ѕ�\�[ɳVЖ���,ƭ�����>�G@:)��9>��9�[�HHĵ�I�(�-��h��$����@����*��b�Rf���>���O�j�Suό丵�F��0�u8�v҄o���ZI]aj�	�<�Yb�w������3�߯6E�hw�a�5�%1*����2֞���,��BΚ
����Drxv;�����?rmy��L۲[�Ϥ:��=��6Yp��j�}5�y}v���C_���x�c�9[>߱���0Z˅ڠh���k2����zqGDx���W7��,�nd�D���{w�b/�^�"�487묰�{֭�&�M�w��w,`�
*��8X�]�{3I�N��j�ǐ��N�٬h���K^�Xז���-��,sE��W^��"�M��+����R��?z��=}�R�*�p��2��j߄�)
M�u�k4ez��9
���7T���S����CaJD�tRxN��:%���La�&��%�����ީv�	^��'��`&>Qe��H�,'6䄷�=��H��1l�(�!�M�^�]�����)vd�Srb_E'E��q�\`����#1J>�� �����페J��U���z8�� ��uO����y΄1+\����'��2�w��k��h$b�_�F5 Jr�p�w�-��x���0;_�V��Fm|�@k�n�gg���%��BEH���|���j�ArVXzqz���tY }��8_��Y:f��U�CQ�t���ѵ��V��a�1*TZNH��GV�����:Ո,Fc7$j1@h}q�^3�����q�h������J�6<"�C]K Ѝ^J��}q�$��6C4��H�ay��tcW8�g�xR��a���p���F<���v ��{[������Ѽ�8]v���z��w�u�Z�����֘�?��u&�p uy�^�F���l�{�K۪��U�V>�u��g�������	��]��4v[݅@d������>�uvi�_���섡(O��<�#�	Rp���Ld�N�V&ښ�b�@��75���D=��`�Dt���i�i��\C�6y ���$P:������>�y!/ʸ��C����Gc�P}9���.`ɯrT�{��E@Z��k�d>nc2�-h�jh�Xh��M8G�\�,K��y{���0"�!4K�~��u29��XS��/G���1B��+��z��[�H�L"�St	v�L����@����B�}������j�$���zC�d�RJ��:^{P��0����A0�R��mG`0,����<�lk}j��*�0s�3�^2�~�h*;'�en��an�P�����%����g��/�S�K�y��Eɱ�_So���/�;��Ǧi���W�bIc ��	��Žxx\����t_��}�U��^�E��tE��7��*�J��j>ظy;�\~�P�V���l�o�t�1Iߘ/��{:6�#.��Qk��D�˰�dRl��_u�{���?�.����4�7T&(�F�_!�6ܭ�̏���E������]�B C�xZ�7[�Ȱ�"���/rQ�0���r� !��>�T)!.�u:�`���F�J#�����t����[��dǆ62��_$4�)F{�WL��x��
��fp�)�h���p�%�e��S:D�w7�3S�M ������"�1����š�)�0�j�6�%���U�I�������-��g�#a��P�ګ����*�4h�b��|͓2�:�9�1�Af?��,q�.|�m�/���F�rDnX��^H�1��TP�Z�����{�ƚjb��ۜ��"�xS�Y+�?n�{��3ވ�r/T��Itd��8�1�(c�v��n��6�Qp�؞$�m�~j%�2Y"x�Н0e�и�[C��(=�/.�� �^�[u�:��E	\�|����c>��b����(�lP֎�e��P��6�=]���e��ն�M���FW���a��vR.�J��N~:,�Ci0�V�$�����/�Ȧ��¨��(V2��Чb���q�I�_z�ɖF�Z���e[��+1��7�$�UeA�
��D��1A,	�:��	?n<�#���=�r(�e���mC�-�U�����ko00�:�f�������@|�=�kJ�G�D1�Y�<Qv�$�Õ`�#�1}�y�p�_Ru���݇�j�/�(?U]p�u9Z��m��0^MŘWB[�N9�W���ddwr�����Õ�ٝ!��'�^��q��kH/H�ɽ�}wT��'w��܊,��m�v �wo�9)��"���Y���hSB#">t�ݢ�t�d�b�3�������gC��zq(f�s�!�iX�}s��V>������@����f ϯ����E�}]�H.�[�r��8�^% �yK�̜ZĠ�6d�m�Vu�D6�Q}�q�z��R^> u��7ɕ�GI~Q���q�Z� �ǥw�ijF�"����o��7Ҏp�(��1�|��� N�>�r��_Ra�,
�_!��P�U�_�;Ei�/��G\e������D7%M�;<k�L(^�I���ޗQ�����~�\2�EmLi�;��j/#���?8Ù@@���n����2����mߔ�E��rh��kB+r�v���f(#��<�}��H�n&�e#mXX_Gr�	�[������#�M�g	pr�$[˸$r)EU�_
��d��|�T-0��2���ڋ�s\�ٝ(�x��f� �&;)��;6*wh"t��:����;T3g���"���&whha�a��4�T�J��,	���b	6�=�`������<�J��kх���m� jd�n� (�!~r��]6.F1��*Ґ���F��/��A��pX���.�p�M�7	$jK�R�@W�u���r��!�*Q��9�pFB&�S�GX��O�Ҳ������qj� �#P!j����v谬��g7�1��n��K]\��P%�R�����������g�acž5G�%���I��y\�ÎoM.���iT# ���׍����+Ad�|-�.h��{(��W����}ƛ ��Z �{���X+h�m`)����fc5?(9�0�.Vn�����\��T*�����J��kRQ�$rK�h���6B)O�g��#ɷ[~�y��Q -���ȹ�'8�z�uY�dd���� �e���7�M�	�߶��)�v"��fT����;�[K�z�J[4PM��Y �a���,��:�7������ye�!7�����P�oet(�$ϯ���:�`
h˘B����:�D搃%tY¬�H3ԝx�|�8�±?5͜����L�B�w��<��]9��4ќ�Y�U�ũ��mE�]���<�O��;,O�%���|�L]E�I��%|��>i�S��	մ�sPP��{�ç�������9�v/��Y�,t�LD'˳}}���2)�^������`o����5DE�#��	��KQ~g$��"�n�}���-"CD[SW:�:Eܪ1�r��G�Y��/XM�4d�w 3�
�������}R��Ͻ. 
����?k$����{�9@D1U�_�Q��-����0i���^^ʑSd����#]�\/<E)�,�m���2���虗-�g�G����'cm �Q�g��`�xDt���w�Eڙ��C���-����_��;����rK)�!���M��dq8!M�+C/����E��©l!�D<M�?�����3<�״�����1q���X�+
/rj��E֦Hu~���Lm2���I�;K��H�Gj&��zAC *R�u�<��q{�Ÿ�X�E�hj����6�Ԟo�K3�m�����;�2�U�΅aDǥGԮ����W{#dp��"�~��vm�W��	4`�5��(��G�A�:%~�[vl^��e@z�3|ǬNC���b� NX1*I�w(�odD�lh�'�@���$�%�MAB�&���U��?�Y�R橒�`��9�k�M�+�4H��i�������u�|w���_�����G�y9Ͷ#��y��a�����@��*%\�q��f�(��#��dO�*�W��Ӕ� �Z���֘�{��9cc�X���<�O�LI(#ۡMN���%Y�x�$�0��n�]�/B'�ZN��s���;�T���쐩۷\ ����m>2�c9=B><��N��e�l�b� ��o.#&�<��,�_�Bd���vH17�'��܇��A�y4Z��A��m�=�7c�d���j/~���.zj���Zy��I���xH��J�5��^�gtp��wн����fZ'�l"8�,�G�'P����	���8�q�mz��%}��1"��?ç��9![]���X<[��NY�ět^��b�pQ���h��%�2���?֚xh��@����#Q�&����� �3Z�D�i)��L=�#�gM�*�Y�dg��h[� �!�\vK�	L3ȁwɥ[�@��]��<L1�,��l�'�<;Ik�������OYN��v��:UM��=��PY$�W���A�[b��[�Kr���5jm�K(SV�G�g��ߐ���\�WC�XK�$�^� dS����|܁�uL	I�u&
6��Dr����*��{:�D����ZGT��C�ѵwbVl���}G<$�i�|dE2�F��W�5"{�/�">wsR�ٍu��q�g �F�_y���/: ���B��:A����a�I7CK��悡w�O��C������vS���?券�q(EP��nȵ� ��`�,ط(:9)�A# 8�0�'h�:0�/�GV�uc�� ��K�k��+5�$��'y�ap�=��v ��ot)��r��s����1����y?�K���m��)x#ۜ%�� (y���NvQ�=���Iq��Ii?���Du��uiϦ�ŧ��� PFƾ�v=��#a:�� Wº�I���	>:�1��5y��N$ai3oY���hQ+Ȉ<�`�_���JE��*�{d�����mT�$Y߾��>H����E�������԰+�j~'�4~L�5�rO@*�mb85
ٺn@�9��)�1f���h O���ͩ|��-K�4t �|���[�uK�EzyT����k��x���/N=:>aH��^еXYT
vS�Q�����fιcL�PO�4{�^j����
UO`��r�~~D�|��%�5����p#�����d���������E�Pw۟ʎ�E����<O��]�g�wP��ֲ�u�%�˔2�N/�&|��:�}�2�}q��� ���9���,=��lxLԃb~%F(�dD8���� �I�f)
 ����$���	��P3Rz��%��#7o�[n� �bz��/Jn8�-㳿#�aI�L�%O@�����`�~���걥l(�	��{��I�����a����7b�^�
�e�K��%���X�*j�}��<�h9���*_}��0��O"������A:$�����@CX'�IM �^���P�Z�p{�QҤ�� �Ӊ�)�J@<EQ�@��#����^_*�`�e�A�up�h[�h�?	�~�}�
ew*����rm[�m.��.O��efX_n1�2uߔ�A�w0D�%-�/��񕖘��L&P�1�ۧ�j��c�~�Z��Q�U�'�Q��Z�k1�Ƶ�Pz�_�'hӾ_�G����uT�����\OK��{��{bC�~'��3j ��)/��2+ �����K�ж��ǧ�Q'"��}��E;f�C�3V(�������x��D!�]�� <]�ux�80�lv�2�"���Q�F�G��x��Eu�,����y��eY��BrM�O���RCy	�/*6�NB�����鉘�t	N�v�^/�2����X�I���Ы��_�PL�=�X��n�����U�lMj��8M�6���ʑf���{�P�����F�O-�7�P���X�"�x1y��^rh�jon�i��� �J0�_�i���4I�ψ1U�X9�	��:��qPTv".������F�@us���G����55��Y�mx�U����t�[�%��� �5���&U|��o`��
W�V����ba�q��<�44Wc�8�8jҠ�>x�T�M��R������W�@5C���@�I�S����j��9�@���c��r�jpi��N#�Rt���l-�F#�u�g�y�;,�t<�g��!�{�o�c���<�K%g��cޑ(�M��r =�F^����.F���m�_��m ����b����Kؿ�e��>��ϻ��<��ۄ$K�e��9{�b���ٚ�|HPs䓸7��cs/^����iC���k��*}�<(mp��ϊa���������St�l]�r�Rl*�q}��'/�6��136ޚvנ�.��F�Bv9�1��tIX\�F@Xh�4 �C�K�. �L0����<��/Oʗ��8f%BP�k�؁�-�PVI@".&{ھ�fꚟ�:����q��c���,,?#�*bd��a�$�&��p�A�0йv�4����Ԁ���SU ��a d�3���ױݡ	�k�\�����[��\IČN�9[}��[��
��E%ѕ�k��b��5�F�Q�[�IO��C0*�q͝��^ӖJn�s�ee7ʒ�z�ծ�M���S/�G���Ul��Tq�z��Z�H��?Q�Ȕ��C����I��Pة7fg|�N�����&�4�d���-���]U�M���0�G;�1<��(�/x�?j߲�d=��+V�Vۆ>nkְ���^�猛��^[1��~�pJj-�G� ���^�$�o�k�qY��=��g���i�S T6��1P�@IGǠ�\�ӊ�Mg�T--Q����������P�W7�Qӹv�C�����6l���u��㏻X-j5͍����K���_U;��J�����9Q�Y��z0���?Tr��G��]:�MlmJ_�je3v�	��"� ��U���y��s+ȈE�=\IX?�Ba���Q�p��=a#��Ůk�ӽ>)d����8a�c��[�6Vѳ�`���m1-n��U�h2��͂`�J���:�;ic�����!I�e-��y?pp�AC��w��hUA���]x���?���/~\&�ƪ�M����ǹ���_��!m��rp'>��J�o}Y�URq!�H'��ABu���!=j�lm��r��nw�5#�^v{p�%:I3B�T��#���`u����rX������y�/::��ù4Q���}u�O���y�6����CpQ�\���Ȍq����,��V��Ž�e0b�4�鿾��x���g-*�
#���h"9E�x	�D&���hȼb��������Ş�K�ۡ�i�/V�/b��Ä��}�̲���˔����
 QgE
� @{��k�h���Qn�<aΐ�sD�6A��� ʹIN���1���G��[�z)z%*��rۇ���G�^?��+�x��̫����.q]Ȃ BO��B�Ϝ ��y^R��@�c�XU��@���>�Q�U���e�K�
���<6�qB[��]�]�aPg�V��Gd
��ܤ��Y�>�*����]�����	t�!�]W)쌠��|�6-}�%�G��"w�����q� ����ò���
��:Ԭ�X�PC\8�CR8RD���Vy�=��Zr���@<����և/%
���B7BJݳ�Ue]��g�n>T�-��:��@�/U�k�]��g�*��wo=��]�l�v#>F�BE��V�m��m����Q���Q�̺+w��r�ߪ�l���ݳ1D�e�a���z��
�<*����}:5�ǽ�%������dk�*xhB��|*W�y@jk��']�0��/3��ͧ�#lRC1��E�@:o�ߗ�v� ����u ,�1�lų؆�3�&r<�YQE[���\25�c�o�8�bg��1f�
�O+S%xB�W�F�֞,W�9�V���%�S*��d¬��̎�b8����u�=kx:gӿi[�L�,Ղx5iy��x�Bs6�\g37u��EY|^`f%��u!��ki˟<Н�NX���{W�����;�a����[�)3� ��@���v�(Af<&4Y����o)���O 
<0�]�ɞԼB ��Nje��:�u���
E�j��_28'������ų��e�t�
ի����uK���T@��n�QN41�|�,�� ��*kؘM��rw���u���>H��8җ����{��0���� �|�;����$m�
��2p�ֹ+�_ߝ�M�wYD��~6�)
FX:D�i�J����K�di3��7��[i�G	 Y7�Qh%����&k
I]��=M�%�2��!#�Q�4��zA�>$����7��0�^F{��g�:2��q���*s�@.
��'{l&�b�m���+�>Ɩ`h�	L�Q*$����ށn��G��������^Z��R"q��;p��ڌL�	_���5+�>�UM"�Vȥ{�ߜlԆ1����.�
8�yn+�l�DD 6Ⱥ4�W�	�M���)�_紿�RW��F��凢M�Ξ.l)����t�g1prR����l��xs��ؑN��|����t���T!���U�a쁆���}wd?� N�4�#�)H��˱�Z�XNq���ĶIqX1?5��2�"�Ô9�$�Y3X5�q���=Uo��+�I���OJ�AR���)9c�zS���n�^bޠPf�H�,��IYi�'2���.Wģ�>;mN�n�l�diDC��\�brՂv��8çD��(���dR�n��e@ͼ�)�����ٯ"����q��k������a��5ɡ_��z����hkdc������r��'5-oc��D�V�l��¸��y������,4�j����p����*v�_M�2�ʳ8�b׶�-D�дǪ5����~A�M>�B����绑��t�~����(7��H.!��:��g��U���cY|x�S���[1|����]F�D3�M�=i@8?4])����M�]ߴl:�R��>u[e]9�v�tO�_kg�K#N T�I�D��-������#��#�td�[�r����1��jP��z�j�)�0��Nd��Qh��F����+��~2b�9왧��>�>�eU��P]Ə�%Z2@�![���`�\�[aj9
]MS��)��Ogq�	�[a�a@�9j����N���a�)`-�S���%�I��
�V?�6r!a[脮�j@�c+��G\<Y���3f��E��1�>\nD	�[.�@���3Aå���E>dU��'�i�r�	��K��\�}Ċ��w������p��]�����D�^#>l��0��'JcCҔ�<b�BѰ.E������i�]� �ӄpY���:*OZc`j��`"el�L�ˠHs �c�K��s �/�U��t k{�?�ϰ�$���ئ��R8���8��m)c�&�ή�$�W�-%�P�E�%jp>�ba�� Ȳok���đ9�Z������di������Z���K����}_�DU�[�x()i�j��o"��� Ь-���Z�n�A<�n��|E����Ń��uή,clg��,'#��ڤ�z��0nG��jE�mʭ zK��Y@Wb{���*t�N��j�q��q�p��y�����W<6(?��^�C���g�k�>9#�Q:��s����,���=L*���+�v���I��gPR���u;�x.�n\?0�*e��#�fs.��d��p��;.�Q�c�=��Y3̿�6��	g��^�丵wqp�<
��ٱ�c��~a��k���=+��{�ʧh$@Kq��t��/4���/�L�ڋ�����mB���fMr�3�d���V�nŘ���F��`�2Q��� �6V'P�&�1�;S3gF���+�����:.��۠�ed|���*H��^w.������S��55���{;��+^�Yv�{�6�E{������s�M�87��5Bʫ�&F�}�l3�_D�U��]}���6�븙�t@gp(�_9frh]���_۳2ڶ'B�Zb����vC�]�g��f��Jw�l뾎�#0�j�F��*c���d?�؂�xTf2�5����Mݒ�Ē�����7�.pU��ca��G透>չ�U�Q>�P[�ɺ�b㓜���⧫����'A)� 9+����x�7뷗�u�i�y
C��Z�#�2O%��hy��0xY�6��UKPڴ�t;��\;_�36����j+6re&���%�z����g��Ex��[��<�� ����`�'x暱�I�j�q�O�,�/��d�2@��-V�y��&�����qz�A�"o�Vʊ�(���sK>[�-�F�e��埾�n��SϏd�'��PLs����b4 Ұ�qx$eWIs�f�`#^�H�$�w�k
��m��3?hf�!r<�����ؿ�������vA˦, �]nA�A~�*�җp�"`22�:9)�i�~��$�a��*���h����>�^*G�d�leҊ��P�%�����+{�ߊ?w�B�M)m1sm�G��䝩�.�������w�����QʏK�����B�:͗b���^��q+�R�b��AT���G�_Q���$�y?[s�A>w���Z5��M7�.m`?�ыg��Oz��Q��F>Ca��L]�������+�ҕ��r���,:��EL��lI%)��3�ۡ�31wYe���<�P@�5�&�&��D��5�K�[��Jz����A_���z���1Y*�A�^���Mv��&n|���]�,��=d���:J�,�ݬ�Ӗs{g�C4����!$�|Zbz�iNPZ�W��Y@D�]��:���f��<�>��"M��@�r������X�u��awpI�;8`�C���z�9Qs�l�����T%�Gޙ�K������Ҋ���M��3�T����]!H)eP�����v<�d �&1l�";�&'�����m��(�f1~��f	��Gp.��y�J��2
b(�>��N���PN�?������c
�o�A��k`5B����N�X��JIQ��r�S �v��86�
��ě5�si�f�m���}\Y�&F2A\<���v�V�f*��K��<�����&�CX&;J�g��D���aM'���$�p�l�}L�p�.�x�Dvm�,�0 �&��x]E}��_&������gV�x�9�uR&#-�SQe�f7�_dJ|�YL�3 �L����3��W�ٔ4p���- sot�+e~��q�4��Ưܹ9ǿ��:Y}N
:Vx��yݚ��1����͌.�F�P+F���9 ]�'�̔Oȳ����^�ڈ0\h�z6��E)����Q@�c��ν&���Dj��f2NhhX�;p���Eb]�1��wF�g�	,O�b�fdp�'�*���_�[^�?w�6wzr2�~\�v����d@`��:�I	�`R�i�el�X���������~� ���BޝZ`[�8ۗ�u:Zn��"u�O��0fL��Nީ����/ד�"��d7��Z�<El�n �;�T��imq<��U��~bR�]�%�y�t[����׶��/��b��J���@w�����<?�gH{���+�u77�](�0L.���o�n��6 ���#����4ajU���G$��,��ưtk1k�5z١��:=���C���Pz�V�#XW�©�{�6?2|Ӻ��2R=�Z���ؖ��\UIQ��Cl}'6��8]Y�h���RM~�t�3s��Tݸ%8)����,B5<PQL	��eduE �;�7IZ�[��#i��_rמ?|�/�u��"+T�F�ѰG��߉7��YJa�4�O�����gcT��C �q��-���kd=`�u�t�6B��3z@X	ጉ�~�8	�R9?�C�Z�s�k;�:)��`���n���+W)���PM�$Չ:���N���h6SD�������*k3}��\�Y�ã5,x�h�(��A|?��?���B����B���i�1>ٯ��	�C���r0o���ȕ�:��P��iu�U�L��p�
��u�~\N%s`H���L�}��B��;PCIdj��G2�XOmo� ��3�E��B>�|ҡ���M�g ㇽ�i�KIc��3	��]}.���i�toԎ?Ħ\����0I�EJ�ƶ�B�Iڳ%anQ��؁�-��K���ݐ��F����SP��<��W��g�����)b�?��1��T���*YV=����&P4�.Ǜ�=y�^�԰�Jރ�qk��8�LwE�����e@�����_�7��29��,ַ�H^�J�c�����TS��<�C��a?i9S�=�OļÉ�_�RK�ka�(����
���ĸ��H~��ψ�>��8{Xl���kW���B�>�?L�k�{�Tp�c�
@A���*��6��&�������Mzk���.3�`�(
�'�d�~�㽇ɘ�,��T���A,��4�G��D)g��_�XrR��ڵ	�\��"*�k��sl�v�9e:k�Ne�!]�L5=�L>���x�B�xJ-f�.]&4-�D�rj�<������Ȏ�\t'� o��f��

Qt�9��]�f����Y��ӝ�]?�Hi��3I�m۬��5MN�7~J�ODD1߁�ΣR�#�+w��7�"��5d�k�.aἤ�3���.,D�%5���T�LBLp�щk�NR�c�V�>�����~�Q3S��Zq���ҡ�ڟ?w���/J���k+`w��G�0:/�iR1��ps2�짭8����&Rp"�0�"�ۢ��;H�a?��ub�41��)�G3}����]lVy
���l��n�v5#��'W\QC��I0�K`y��@��"�콴H��_���)W�1���]����fvo��qz��C��%s+�p�������$?���Y��^A/u-ALb�����CuXV�F*�)�R������8))Z��92�j���t�"�����#+�`�����W-������8�~�
ջ�Bg�2��mc���5�Ѳ��lT�OOoT%p���	/���mvPO?i(����(ct���F����_��$���b )-�@C�}̪��z6�z���,����!$M�G<�R�q�؍j��;���\�M�X�J��8�j�Qm�k��� $3w����uU���	��!���]�֮�tk���W�t���̮\U�8�R����ٶiP���b�YK�O�d���˕`��\��,������*PVǞ�
�,�D`�����\̓~t'��y$i�Pk���z ��9<��ů
�;�<�P�"�*�D����dg�0��hD)����I��EbKXY[���
_F*���c��j��n��@� �@Q�@��=��DL�X�p�?�W���]��* ��ڝ�b�����w_m�T|��Dn(`6;GLS�ƀ���%���J��Á#� �.��8�7g_������?���S��*�	�39��*R�~f~�_������_�(옊���z�e5��z���qED�L>��1JjǢ��E��D�'b/�5��Y�~��0�����h܎Ti�&q=�R��Kܜ�xī���W������L�����3T,�;�1b\U��ը�y�`�TR�����R�Xp7U��}
RX�y	��aE�*���|$wc!��$<��ye���̕���+��,: ���>���`LP���m��#��3�@�|MgTgF�슦����8�3�j�H�9Wթp�6fG�y�V�C.!J��F��s)����w�a>3�<Gdc����ڰa�;�Z�65l��Sk��ހ�Tَ�	d�f�.���B"��#R��[�c�!��`%Ί���h���*�q(�+Y��M���>�I%��Fq�˸_c	F�xe��M��R�[k�e���BQBHtۺM:���Ƌ7��!�6�gE���?m@�#���'0���7�d�5G?���P������ńOz2���YݫyϬ+̔I�b��4I6?|̷,I|^�b҂�U�,�^��Ź@��v��ۆ`88��	vb��Q#mr�J݃煲|��	����q�9ˀ���1�|�]�ބ=�[N�e����.<N
Z���A��с۲��\8n�o_p7�ș�mN��v���9h	\X{�EL`���3��o4�f���!����PlD{�
Ժ��j��ջj�|k���O�ĥdn�|���I��s�  ��X)��6G��Ė�3r�e@w� )���"^���P{�Ydh�nx�0b�ė��=¡���>G�
"b�xġ�"(��?�o�i؉㯙f��Տg�昿^��e�8�7D���{FMb�yZ@���+�g�9��f�J�C�������/� ��������`����}�݋.�2ȳE�J�%a��M�b#��^��EP�e�?���b/.d ��K��+ԇ��|1����e��
E(��}ߪ;rviɤ���yQ���%�l�:%��Z�����m�c�0�d��'f��^!���,JP6lZ7��@:�u�^���<�Ĵ���_`ܶ��t��&�RA��r4���;c�#�~_��Xt	�`�OBM���iB�]-	�t���5:j7��M�#K�����̗g�R_���\���y��{��D#`�=Pݦ�.�_�C���"�	N��=�%U��r�r�>Zbu�@���`���Ģ�w���r�)Eq+��yi��(�Ƅ��ǭ���f����|o��$��Q��#��a�^��Ս�!��q���3�-a���X#ԑ}ު��WE�������G��X��O�pҠuG�� ���i��x���Q�2^�����?xF�6���3�v��*<�ߨ���P!W۰"B��WL�ͽ3fд?��3�|xz��OX������&���s*�k�ut�77ȧ�r�a�MوȾ��3uv�:O�ـ�3�-�� �In���O��.��ppb⢌vSy� .I
~���"��#?y
�1��3�>�̎��=O� ���t�$�r|p�1�!�&v��������a9J��g�������� G�(��u=pu� ��c �:�s�Қ��,.����s��Қ�O��,H`3K�G��!>��1Ҥ�YK������"R��y���N�vL2/���1�)zM���^����H���sr}�;$�;#L�̎��}�"s&�OQ6)���/RFPC�mmE6	��w�����c�$����v�э�WM � %�P��_:o��`7��'F���A�Վ#���lud��_�l�򭼎���7�g��*��������]2NR�M�\�#*��ڸ��{�k���vn�Ƅ�eم�'w?���G("U�Ɩ(zy�W��Ri��'�Hx
���==Do��Eu�/}|�;a�Z�t냮�� XG6OYV��*���v�������=���^BJhF{�i��a����y�����$�'����W8B�F��S]����n���֨�-��2*����h���9^E�m"���h�$��	Y9F���1Q.��T�=s�@������o���%TB�U���r{P�p}������;
��)�d���@�+��\U���C�bM�c0Z�M�Vt���H�@�C^��1�7 i{A�� �;��j"�xm�f�x{V�f���������ƕ�5�T��^�R��8!ڍ���F�]��s ]+v��(��2 č����Ш��+��[ƙl��zh&�𹙗{�����O��?|6ާ%<^��s�`��̖�l���I:g������-�	PU�b6?�#�;/��?=��C_��q�t$+��}̀7]�C{����<oA��&o��HZ��5�P;�0oZV[�l���Z��ӓm�V�'%��lK� �$� 8T����X�@�u8�( Lcޖ�R�t�(?3��4���C0D��R��$�F�B�:�G�*p�M�.h^%��F;��C:���aiIB�ֶ�J=�x�)�R8D���>�nt�|z]#XHwsD�_���`H]���ķ"%��5�AD]咀Z�]f�cCH���s��F'�W��aJ���zC
r8�V�jF��DjQ������=�U��?x�#�{��S�����?&���L�����2���r���}�h��;�ˌl��%��*i�m�����)��J�)b�aаǍgw[��
��t-%x�mN�# :�գt��xC{e=j8FQd-�	pTȵViؑr��Edi [�0�B,���d�;J��a��rWId�ҁ����14�w@b���wi�R�1G��Е��F[��i9����S�0�z�0~�8Kk�ؘ0)����tIr��~���}���a[����l<�,�i}Q��`U�7�x@���9�AW�����6����ոC-��.��=f;��FgX)��e�ڻ|W.��}�7p&�$r�m�
X?h�!��&	��ȭR�.|�9Gߓ8��kH�$H���uS��֑�7 ��1��2àX3�K�����C���X��AL$ri�M�C����-w���yGW;j��t����es�	:I��䳠�3��Y`s���^�3��p_4��(�����Xz�k�7��j�4���]s�R4��[j񮷈,�����(��WL�}_V������I;I�3���CM�O��E9i�4���&P�x��F�/��$�����ȃ��둱D�}�NMd��.�<+�C#i��P*��sG� ���ҋ����cF����M�}=��Y����*�J�G$�?ew��P p����ũ�4�R3��h{<<� o�+�����T�G7�X���E�]Y7n�Gu��֌��Z��/� �m5;�G�uV�^�S�����0O����Bv���f,g��G{��0<�g�^NՄ�ѥe���sO'#� 4�{0�X�v�5�'�_hk�X��WY�rwn�Nn��L��
c�ȇ\k�I�uv�����Ʒ6>>���&!"�F}}ɍZ� 8���lz7��`�Q3^ 7F��m!yy!-O딅b����#�9�*M?�Aꑄږs����UKm��A1)�8�y%m�۞рB���J�a�$��� H#7�|,�Ľ%ֺ���BL��ϋJ��$����4��������C�1E���!����>��囌[7�׺�1��5H�k�38�%+�X�$Khe-V&���6��ĚuT�wJ8�v�_G�P�΄�ə,��#^]�/�sM�y��6ܹ5tz��b�ϧL�A(V^�4��6]��B��). /)�<�yg�}�z���
�5J|G�/��AZ�5�.�7�������' �
C,,Z;��!N��p`��dX�Oh!`.s8L���u��1�z��T	>ܡ�*��	
�&\��S��[\�}S*�����[�����O��}�n���%�Ο��Z�G�{�\����B�>��o�����6m6�.���KW�@S�|�$%�=g�v�qy��>]���kac�BS����ھ��g9�W#*j�mpWHQ^�10�]٫o�����ء��a�rk�]��h�98!�o8%����Q?�ˣKbM(���9g��*����*�n��t�'Yͣ���`e2<�mj���E,b����o9�"?�j�R�s��֙�&���+ʀ����#Q ����vq��Ǚ�r�,��r��&���k���(8$���� �������DY�%�(�
|i4��!�����ɹo������ik� ͦ��	Y]f�X���_��L�D�j�Yc�疧݁Fט�	R?��mQl=�v�-���|j��`G0��j[�%2R�KzTqx�H�};l����}Uj4^&�W$�(�����MM�h)N�g�M�p��ە!$iMm�i���L�>h�to3�9�O}L�#ᯭԳ��$�L���*�$<t�6�v���8'*�& t�����{E9�7@r~`�^cW.�'
'4�H͋�,<BZL����-����ge��'<����<p�OZe��}�Fx�wf�\�)���<� (�'�D�5�w`d�x����78��=L���h���)?F���G�"�.�Y؁c�&�j��xV��VX���9��s�@������?e��_���d��������Rd���Yx���mMI�]X��(��x�@�;�Ս��*0��:��� ��ì��9k�t2tQ����D���N+���}��e��k���aW����pӌfڶ�3� Da�T�@��V������ŗ�	~@=�(#-~�j%�Q�������:i�n�g��};�BBa�ū��]�p5��O<guRm2�1b5�q�����"��)�0�Q}~経�h(�Yro�� ���҉���:�U]�teݳl��?ީ���s6��P:J�\�T� �7�P�I��<� T,+דmW� �������jR�KK&��i��kK;NLJ@�yv�A��?3���jd�������Ee�F��*���9���l�Q��r�
�;rEb��VF�0�}'$��c�װ`_(=7��Ck�]N7���3��}�\3*P�J9����bH*����S�f�븜[EB�+3���7����=�˅ t���r)J���hy�5z�zŲ�*�|��Y�_��r�_�hB\�<��n��Y $�!�AkZ*W���Q�������=�=lr�� �@)b-�|R�0��0��q�I�@�TB�Ў��b6攟�:}A"_��ڤ�����6>����L��	YV��?�Zt�<USC��t����WY�\�+�!T{��� |���0w֏BC�?���
�%��߱!�U瀳@t�4�X7��K�"�0��������[�j�F2�H&v����W}�y��	l>��>���t��$Hp�2��O~���\��as:������!��테��+JMJj��ʮ��2��?�*�������� k���̟0nǌ]O/@��bvO��T��d���g���,�����8pv�5}�]��dD�{EO����	�Mi<�̜�����֚�:�DE��ʍg)kIoT��r��������"�L�Θ"od^�T�Z��%�$�yy]��U����asJdY��D����:!��������y&��B�������.��=�ĤΨz��f��8�6�0ג��C�Z9�e|��ȱk�Y��|ᠯ?	��EZ�l�v|��F.��^�w����H3b��G�[ߙ�զ{ě��n3���ñ�BI|$t�j�����a
�p�qLz?��b�v)��k��Se��Љ�h�g>��P�����;�}li[<� �^�<���䮡��Z�>�����T'��_2������^��)�����4��7�� ����p�nD�k�PH�Rj	�I*�]�?P��ɰ�������[KD������;�$<R��Of���,�d.�Ƭ�\5,����
�w��TDU-�]^Ț�{Ա<E�19�
�S�;��۩�,B�0��>r2ej���8�)�*?#*TA�����ߝ�����Y�ã�^�ı�""��pU�K����B#��̻��g��r޲�T�N����V���I�0�MP^� cC\�>sm�箧����a�u��)�jD�>wS�nL0'��;#iHp�(���M�ܩ�)�!р��'>����$�:^>$\�����G\� ���d�Z��g�Ǹ�ع���n6P�	eb1k5� ��
Ƃ��g�T����1� �M��Ң^
���ETz��V��~n"���ɱ�ӟ�*�uy��I�蘋��&W�{R� �/�Y?r`|[:��wϤ���|[c{�P'�a;9}�k�n0���T@fĨ��N��nsqA��%��=��	9�)�P+:�ס����O�1&�D
��GVªVA���-�4C����"�����u���앃��i��l@�&��bo�hEB£��e��䵔�8�V�T��Uџ�	���˨�`w��t#�+����*�	�==�z_�{�.��H���C����Nk%#��mn�RK_{&&�����Z�7�Q˘)7�.R�	7|��o���x��̖֕I<�z�&f|�@���h�|�s,Bt�s�,^�cnoTjD��D`�o uh �KɉT�e��Ta�\s���� �F�?�PCʗ�$���'��G$:X�:֜yW	���s;�ȉ��Q�8�i=�~��ً�VH�m��7���-�?���X#��_o�ыeW��4U�c�

t�z�4<�>}����Q�ي��BC�E�`��!��C�ZI�%1�y?�e7�"�C�b	���8K���O�A~,��˛���U6���Q�/�4�8���-��\e��7ĭ�Â��kb�ƓR:_���#n�8,D!�c�k÷�#�����`k܅���}yF8�>/�xL4g't�l:��c�� 3���4��fE�Y��3'�p��2�ˢ��\G�X��íuW�y`C�CV|���n~*��x�אֆ���B�8�}�;�2])8G��u�I��[r<�ъ���&3��WFD.zZM�fe�iOyo�׀9�� �l����5s�4�OC�a�w �J&ļ/[�;����S��˴���t.�L{u�#�B+=���(\ڝ�-�JJ��Wb5�����Ꙅ��s"@r��n,�h����С���o��bY@eM����ָ+��
�p����|֢��tK����'f�?��fp���ċ��B�U1�,Y���ͥ#cXޘN/�>��kO�7��E�3�����6yX�i?���Y(h�x�n���J��e*��}�sL�m�6�&�h�!(�0\�|쐰N���>3a�-.�UL�gNc'q�'C�^l������J�C���`�:���g��Nk*���^K�M��^_���-Ny��y2�ss|����(���#8��O�B�2p�LSu�E����Ϩ�i8�����E��^�b���6�@��T�>Q6���ެzӫ�s�� z����&"I;)�!�"9{?e M��''�Ay�Hp�,�
�����Ȣ|# ��VPwԹ�OF�@������;�Eԥ��SGԼ-]�[���F�d/��}�����@[L̩������w�ƴ8ټ��3��k
��'�!�Y�1
4����#_��g�x���-1�[�\�ޏ	���NW��^����!&jOSK�.Ƣ�xDP̵vXq-�I�(}�\i�i7Ҋ!8F��jE��՗������YJ�p�3�:��VO�bt9�	���)�X��B�Ĵ���d��d�냎6M��8�BHD��/�k�s�_0b��z5��Lh�^i����9�����0Cb��[h}�RYdgM^��#��8��r� �`!3p����oe0b��F?�9XЪ�,1���j��:jOJ�\��5��2�[#�J��#l(�!��r��
g��E���,0p���G��bTv��G�Ψ��B!��+L�~�Z%�N�����$����,E���g�Z �aߤ�`
>�M
���%��N��Q��J�X��[�!WE:��W%�.���r�7w��2�DP:�g^;�^ET��I`:Pڶ˷f��� *\dȮs�K��P.b:��
�PIhe�t7�ݛ��735�����҈�����p,B1L��~@yV���f�n�W�sR�bW'KǪ�NZ9�u��T��E�X��)o�6I1A|�?q��X�r@Z�>꒴�t%�'�(O�Ǵ <��:i,%�n�f3��Q�,�Q�i���e}]��wO�(�hX��g%tL��t2p+.��='
��M��8�Pp@B�Lv3�`X]^�Ck~�J���t ��G#r%�(���V��F��ey���Oa��P���(�
%c� *����&;��x�F���+��t�Mu�(Л��Y��׹���.�;�����t��n�!p�I��egHyX�e͏U��H2w�R,�A�71�>E�� 'dݥ�Qϧk|��^	�?ra�����x3�? �q�­g
=�`��pשt���������w�m,+�oj���������' =7[.
�NW�$�*Bh��UCqw^�����5���L������;�5>��g�0�5ak��V�6o��K�� b�o�K��I�uK9Hq��t0��Q���u��R++�x��UHV�Ur�V{2��������=��p��-����'�&�A���ʩ�A-iK�RrI����wx��՟���ܶ�����/�9�b[�4E��D�W�_$��f�j�4;�s����3Qgݫ���uz�uv걜6-��ؕ����0��5m|�J�sgpvHhp^Z &�}�+9�j�����FR�U�F+HH���:��tms�ܓ/�s�f����t���;������ʎ������j���c�[�C���b��vmH,.	?u��C�lsiP�Tʆ�.d��pﱳd��M��C��РF>
@�!E��	�!g�_�Ա���� :�z?�<[�Îd��7�/�S���C�-[c��-=��9�	?�g�!G�=ݴ���41�y�o��:�h���)1H�.�`os���N�zyR���`+0��}�T�}vG
�u� ��R�����|(�P��M����KJޜ�m�>�#Y� @t��1$������2����G�\�P���X��$ڄ��P���|�mu(�,Zs:��fhM�Ct_.��i�?���S���c%{�p���k`ӕ��73.*1h@���`�� ���A¼v��|*PF���N�Y"|x=Ϫ���U�9� $F�Q����pn�|~�8ƗF��� ܿ�v^
t:�_*p�� ���.��RΛN�ī��N���+p]>��O=��Y�*�&�MS����B���&���q&�k�7e����.-ƫb$���O~\�B�P'y�oeꖊL��ְ+���,@7-Ѝ(A_�%�Rϖ�T���{^ʢ�?�t�^Ax���8�ը���V��qA	��\���Ka�F�If�����tq�J�Lۇ�9�^���!{�䤌�w5��0w��ϒ%4y֋AY�a���{usaL"�(v��~�Sˡ�ϽT��&�����_N7d�
�4:�~]ۣ�e���L� �t��������3/X�|KEh#k׵_]l��稶˪��)*�����܍K��#h@���8����/4gy~?��o�Dku�v�����zi��2�3"��P�[iB
����nDuÁ�2j�hb;�~�F/N���K�uW��i�J�.����Oz�&��"u����P愕�d��ź�~_qB�?���M���q	�1�⿚�z�+2����c|�QY!�n(�d�O�̨�07Z �j5�?�C7ſϜ&�+5�&fd���f0pO0�3�}�ѫ� �D�?���W��A#J���&?�l ~����i]u��#������{��A���Z�$��O����}��`&ؿA�3YK���e�=��܈��?vY׏i�d�)鶸^��g����#~|�����kiz�JJ��B�D�Z�z��ʶ+���Q��^� ��F��q,�^�JBj�E&y੖��
d�Ɂ�97m�/��;T�r�Ж�T#��-��7��B"�ۊ2{�N��w�n����=%͔���b?��t��x����y��9��t�r�?\z��������Q���o���z����z�Vŝ��y`���-R�b��r"���7��M\������b�r�@"k�&�i4���:�� Zޓ]=iNft�؄D$�ȳM�d�l���oN"!�K�9��W�Ȕ��DC�u)gU~FD���e�4G��..�?�{'��D���8
��|��u�ǯ�9��9#Y�)i����9@�$\:a��|1�2&<B�C���r#˨��d�b�������אe��е�]YN�z�T[ke�8�5܈������S�g��1�j��m�z��@����ǰ�R8��*L�`K�RM9~?t���V�(��yT�:���~q���a���	"#�q67� !�j�7P��r�Z����1=RPfM�wy�Rq@Ā���S���%)�0sf��P�� �������j�������.�sRΨ���>m��VnG���,���N+�n��s�H�R�,������#�z5��
h���._�s��G@&m��&++�X�x�f@�[���f�l�ڈK��1A�(��<Q���сf3���K{�����N?
Ѫd��Ãd�ܗc���g*�F��mZQ倵�Χ#���M�0;�|�]R$�����ϴ6 �-o4���kF�4˯t��]���Lzn�'��b���k�����#�HnrX�3�p�-�wP�0��2yb�L6���aUlA�gL6�<�4hnr*���	XY�L4Ŕ���skywg�-q��Ҳ���|��0ox6�leՕ:y��x'�� W��7�Jߋ	h�N�8��v�w�v"\.Z��u~���g>""���u����U�l�T5���S�@�xC��i�Eiz2�B8]M]G���6%^���Z��b�Fr��f�i[�X:�)�Lq�@���|&ʇA�v����H^BT*� v��fK�'���S!�R����i�&+�sQ�=�*#<ݞ���Y�3�5�/Wq�m9gQ�s~ZcY2%�Tb�����  ��Ձ[��Pl��w�\�')68Ԕ!�Z�
��������\��]���O	/��'R���w���p��9��$�K���p�P�bM�O����z�J�i�s��ת\��������	�F���X"�Q���_`��E�L�x��ӳ�mTBQ�g��5q������B&�;>���J�I@>�1SK넗�9A�������`�"t&�,�Iə�{��g�`v���d���R����2P"����+R�(��!��!���ut-���s��U�ׄ�3A�BD�&s��ލ+�ƌJ|S�f��������{Bldo|�+�t
0��Bs�Y������~�ӥKkz��  �;ZTη/�ϓ���;�R��~=�
R�(��L?|��I�K��������"̬s��˓�������X�9��Ĺ%䋉��Kޅ�*<Q�N�#n)ql��� �ng"���L�o���E�[+�e�I]�^�!�����z�wr\���U�� �Ԥ�'\�p�\S�)��:��5$����<���5��0$�W�����3ɇR&�e�}	�k��9&v�\Y�q����>�B�����
x����@��U��)��%P�\�����H9��8#2�S&MnL�p�����2,�/v&�E2 �#�-���4-��m1_^��1Eܽ.�$@"C����P.�p���p��e� �Se�GPhroH"C�<�__8# .+��ѧѠm{���c+"�I�����QS���������	Ex�r�ݜr�MC8C�B��zoE����Z����Y�B�AP�j��$���1�~e������*A��N�n&s�)r}��$�t.*K���\$g�ԼN}�������ܭ\�Ȁ��g�m�)�B�9�)s�Xk��NǦ24�KCn;+qu���Q�@�N����Τ�ADx�n6 ��H���THw�2a��x�{J>�Ɂ��h�@�_n�J�6k4I��Ue;<��N*��� ����Z��줋==4����VK�x��1�Sw��'��2B j?� �l[��9Joiv��a[n �m���v��6A���.˓�+ۇ!���ora�K�Ͷ?�s��$����H����{���!�*���^�|��״��Ï�H�Lh	=�U�X�L��L��h��s#G�����1�����U��*�T��U��V�$x���d�!��J_�5nb(�����b����פj�T�Fg�Sq\,����s\&�`��<S� <��N�������e��ܢo]�W��s��C����5f��JL��K0 ��;�@zYnQBi�Q�k.�Ù��D/o�����Q>�-KL[�/���ܿ�vG���ѿ�cRRO|�ݙ�X+y�27�uN*^3�Bfӌ%���:�����0u�K�̘��l�K�i\�h\1c�FU
ؙ�.��W�|� ��"��e
���e��d���O���^ ɩv5��:�7�q@{���<st>u�
�^�m��ęN3�'���n4ۀz�VT����J���fv!7 �ީC]�E�_H���yl���0w2��Z�^X�p��X1��S�)�	C�������sM�ш�����0Y5L-�t�������̈��ܯ�kt�EEf:!]WW�l�>�*qn��%Nzh`��ۍ�+��܎���|���=_�������n����rsiCKx���	���T���ن��?�g^�k�1ii�7�{����Z�]!Q��V)�Q�����I��_rdh"��!�nk�v��ճN�,�obc0��3�U�� �ʥ%iJ'o��$��{�|��|A4j�SD#S
�B��M���lbW��Ol�����4������ �FnB��A,�l3=�bA�h�/�z��u.8m�����bmZ�`�h���ty�^��1�01ܭW�!���v�q8}��	����;q�<�k�n���㤅�+�l�;�(�nE�}bVղ_Y
���}t|�������֌�XF�}�.��������H���[�g������}����tA��Xx��=&�P��+�����T����Z���!NP���lJ�(lP(F��W�E��82��
�o�w&��=�Bտ���`�,R¶]���G��1�qs��f�;ٵ�{K3��I�bR�V�6��	fgW[n3����a�4A�\>K�\��D1��97��Ƞ�}zd'�(��t	������>����W�o\��_2���\,Mg�z�#q4���9��QԴ��:��'
'B�a�S�@��i� )�D	��jRh n'�r�N\Ɨ���Ϗ�O���8����p}������6\dX
:?7
��b�Ƿ���?�zT�$��#��<�[t�,R��%@B@�y/��
m��G�<�}r��F�)��l���Uc��z��ƛ�z�LًvE��2�z�"��O�D��I��A%E�Ae^�쮯r����o���ې�X���&�q�ÿ:a��숩^�:O�BMP�q�w@����Bqj�Y��qt)K�<~ Rqx���~�CD��{g��Y<Z�V���©���0�-IS>ϰy�1� ]l�H���K)���˛�'_�ľ�i�n�6�$q<�@�4*j�4R�F�&�$!�"\�؁�������}�d�o8.��1`����EN�M��Z���g*�}��|y��1����\4'�/��:%� ����)�� Ў0�	D&���PE�S��U��o�T��B8eF�v^�i+�`�������&����wD�;狘��=�y�U=1�`�P&����uTW�?l-�4������A�͑Z,��њNOQ��w���*vm\Ȋ�UE��rpf�-L�UJtZOL���	L�yq6��OG��i�3�p�"�؀R�`����� $��dH��y�q'�����o��b�;����F�=ݾ&n�~�^FX�*?PT	/��Ѭ�D�П��z=]���o�M��q�y��)������G#2��������D|����Oj�}�]|���x�ж�}��f��W.�k���߉3:~��\31!+&x��/[a��ZM�P��$��H\�KB�L�dnb���c�0w��}��tm�a� ����9/2�ۨ9Y�vv��֤5�	e ���Qx��]��A�G�Z�l����g�^�T�;8�QG��[AX���֎���n�P��㿛��q��lV_�p�$�^�t9؅����q�óI�9��`���3��� ��H��^�j�lv��jt�l]<$�n���t]�o���ח"�>������%�{qU|��ك~<��gQ��Mc�t�&�����q�XC.�u�{�;��Dc�e��J׹�M�$�MRD���.�dK�m���қ $�e����
�U������ɥ�2�l��9�(@�C��a�����i�5R%a~k�	Vah��Y��".ٳ�O/˂`R���A[M;c���⎜{f7���푉�:�fLYk|-2O|Ľ���sA0�7�6����<,�h
4�.s�J��S���c��U��`�F�i����O���,ٯv����7}t-�Ŀ��8s���d�����G(������F����v?�Iæ�?Qot��2����e���*����H�]a�7S��(XZ�gM��1��#e��T��Z�_����ǵ��ǌ��<L{��~�IT���%^�atvrϲ�[p�3����(7�+qT� ;�A�H�<�]��~}+U���8��wH�X@��njg�fwB�U�ȹs���j�&EM7�	�h�8VX%(m݇��7�;*/���[8�L�! H{��H7]�Ҋ��4_ٰ���ފ�x
T��P�ޛ^�� �����ER�n�@�醝g;��6YΝd��Ӡٝ��V�<L�h�ة�����5Vh-��S���&{��������7��F`�����/�������6���Y�)���[�oG ����7(���C��3gxf�Q�t(!�^;rt��7���+NYbXbU���8��gib���b��KfKk��)v�F��� �	 *�<��8"4H�C���A(*���H=�ؽ���n��=Jg�L�U�^:���R�v���r�)�3\��8��dH�ߓ�
s���@UMZiF(���ږ�齠�v�I}ψ
x>i+D?g��3��DU�o�)v�z�wI"�_�j�X����Z[͔��	�(q���B�&����u)z����
��^P� �i��1��l�!¤���y؎Z8�xNn�Z�J�h�Z�x>�ro윞���^��؀�q�p2ùߒ�Dv�a�L՛][Zx���y� �J5����gj��.�A]���P5���]����9GU��	��i%i4b̚o>�.����4(�2y�B�$�G���B3�qZ��6n�U6u���
�B��7�d�a@���P�\����"D_�����9�3�_�;�=E
GA3���mEr�2<�,
8�J��#���(�8ʷ�Xr���sV;%�D�QGXɥ5��_E��A_�./+�;�?�*��Rk"H���omF&x��j������#C����@wo��7q���k�7���%��2 ���Q�=� ��]��&��Pas��d09�־�|�S���nh��X��������`��9W��H���T�S�,
���8G'�:�qO���^K���m�02���!��Ѱ85>ͩIf�*���w+�Z�=|I.�f�������������lr����:˶�����G���<gS���S�XM�a��3 �O�O2�}hNƟ��L>��L�2���[�A\o�^�V0s{�Zxh,��NX���B���>�9�9��]6ňk�6������[�Ӌ؊a�g��-k��M�JNSFH4װ��K��oO��� 8JB2a��	ex��8�p��A�m ܅��A��b��<���"�~c��L@�qS��l<�G@��v$D�����d9y~��}��q�rHeJ�����M+��������o���&��(gQl���m��F�����WpA|�w�a-#����F�Ӓn<���N��m�c�"�9��:����H#�ޗ�&9�H���vRO8�\�9H[���6��M�@�y#����aS�H`�_�/�GXW�3=�!���zh���kdd��0�h���K̳�Jc)A^�ҋ��;���?ŕS�Q��/XA�݅��J�4}�A�����Q�nM���]�%�Q��3�G{��k��KZA���l1]������͎�
�⢯�4pi��-ŕ�1�ೈ���ݽ-�u�P�v6�|�q�d΢����6��"T�lf�;��]{���؝����E��Z�=h�5|�� 4��=>�Կ*mD��B9��w6�MY�&�}O�p^Ow���	��|�u|f��lM�Mq��(?C<i��GW/z�簸!�)+���1�0��Yȇ�ye���I�T�]Qՠ{Tȉչ�+�8��6"(jYo��:��;�Ǿ	�y�gз�g"�ΰ��gݙk�������rMr�O�f�g#U0E^�D6�~G�OuMɭeE� ,!v�bG9��LJ*��%<US�z�������Y��== j�	����IR�9-N�z�5�Ҿ��	�E;�6cs_~�5"˄�LEF_s����Xˠ�{Y;�@���pH^o� F�Vo���C,��0��Us9���X�V�..��W�>����C�9����m]8���c���T�Duc�R��+!cH)�1Y�&gmƾ�/�N��I1�8�p+>��1*h0>�	���4�:ޒ� |1Q�	)��BH�=�q��4��;�w�(i��mK�ا���^+Nz��-#�6Q�>[m�k8@5�mq���������'S���Y�v�|}LK9z� �W����
yM%�/�l�]���H�ȃ�( ��6��ئ�'x�)j��PW%g�%�9�G�ڈ��І!Q�<z�q�l����>>O$�oZ�-�<����$���hq�B�BW�����`�D8�4�"(�1w��'�ѹ�����,_��E�%gB;�\'�zXw�kDk3�~�>�[%���C�EQy
	�-+�7`�+�Rf��5ۏ>	��k�4�ɗ�4+��cxM�I�S4QfL�j����qF��K�a�tI���G���T/^Qd��j��H������UR��Z��CU�-��w�"�$��#�]�?��|	�aL����Y�#ˣ{*,��5����^)��i��|Z�)�Y��s����v��m�@���n��2B.+�w�g���8{p ��J�D��
�YB�	,2�]r����P"]�eoc>r�1z�q6[(Z'��mbu����C�@��G�D�� \�eC�a@����V}s->_�|*<����h��
����0���	�YE^8�Q��H����I�Ј�B1N�Un�䑒�12B��ߧ�"�7�o��3v�!���<��LH��+�=�ϥC�k��5�9sMQ˚c�w�"����/�8`攈��f;���J�?��Vܠ,�.�ɑ1V��T��IQ����}<wJ�����"��y��CY���[`i@<�M��o��A����J�
�p@�F>�Y��|�v�3#�t�$,��7��nG0��S�-\UA΃~Q���x4f�U��.J].�.Bi�3���$D��O��*������H�A�W�x�����O.L\	S�'c�E!�T�nI��T���2|�qʥ;�$��S��S��у�P5j�����$�s=Y�[`r�����5J�N����j+:�D��qL��w�$����=�>��7�2��"���"�$N,>��PVi� ��^U�n��?�!����񦀤}�0p�����G|>��yI/�e#��G��ѩ�+�]�έ����V.tS���ܿ����8�:<� ������9�e�^ ��~��R+�4'�z����b�i<���h0�vw?�j�5�^�'�P&�S˓wu��oq�+،8�����r/j,�	%Ǘ�P���e����̓��hÑ���|���Y�FF���b��V֥�k:|(���|��:�fQ��VG}{��j`Ab�!�ۅ��-O1��l[�2��H��LSr�$���j&f�Zr��eN��in�|�+��kI~�L5_�=�v���~1�$�J�+�H�«5x9;ђi�[�^	�S �Uq��.�E5}�t2T���-RO�Lg�;�B��"�ȿU�J�(P��ɩG�Y���>kC_������WyoO��븊a�X��nK�d^�u�,�?��1�-"oNh4���L�69F9�'`�h�.���uL5���,w�kT��R�����p�����Q��i	��"�v�W�]NSAe� ��z+�-���O�m�
r�dB,�WC��C��_���̫��$��%�k�
d���W6��E���5�A+@�b��r��c�%m��=6�h7c	�L:�'���U�S�1K�Us	�\-P�/�Kns��,C���Z[k[�����hI6R�f��fv"2�Y�Sf�YKT^���JBA�wb/e�� ����wJ����Ѓx����i����zЄ�SV��� �$J�H�9J�D�_�]��z�r�i�zH\`>�L.��G�|[iA 7B�H�`����I92O�� �(��?���A2<OGc�e����c��L�3D���b-�W�0#㊰p�2t���*� �hז�>y��j����))�={�'��+ E��8N�Z�6�V}���Z�_+)�_�u�0�V�W�܎���*?�5������
;NR_��3O}�i�Q�I��/�gAF�{߭�7D�Y�A-&O{нB{V�&�������]5�&��!�'*9�v��w<C�#t)���l��*�X���0�������
��g��<ic^ r�`Al�d	`^�����֘�q|1�W����]�e�V�6^����ڱ`�"���Q=�3��z ���?��v�$�ۗ����s��t��	 �X �#Y���	��gmeP����q�_�(�u�.���ţ �b(5�ן@�Ґn>I
�
#�w�66�T�0R	��=N�⏬8�-oi>ë���Z?N�������J�ׄ����ig�Ш��ڕ���3}x8&*���	���l:(�	�'��Lϓ����vd(��O�Y�Tl��hr���=R��s��W�A��<f���'��zS-�,�1��N��O�&}&����� ��[Y=G��<�pP!�S�T>%��o�$���Ʀ5��!Ǒ׻]�	LE(\�����x�"+��>?���:��[���$zg����Tѐ�S�2}1����Y��Y�ݺ������QS|;S;,kg�+z`ՒLf�iu��Z#�	ѥp2f���V�����{CE������T{h��:��s~�y�����d��a��Z����ʴ��u�	��Fj���|4�5Y�T-D��9(���c$��0�"���5.c�N�{ǀP�/Q
W	�-\� �MP.I?ev�
>+#�`��O�Շ�0���`�ڏM��jv^ �&�f��K�����n	&xU���h�ڈ��L�Ch��0�:�Y�H�r6�R��d�;��DWu��������e�������1o&<ڷ�5�_�xXO��g�bx���G�����<:F s����������k�����C�ł�׍�lW�*1�b�Fa�<�L�SO l{��<n�|�B>�i��ړC�O�"%	�K���$��Kp򁖖|���Z��V$��� {̏�&��זӒ�c{<e O�����;�RK��MA
5gb�KV��-�7�]�HĽ���I�
v������������Vi;����H���Q�\0����	��'�����D��L!F�;�j�vg�v�ھ��G��~������t��~Ѻks (30���FDy6�ak��U~=h��ARH��H�Av�=��zC~O�G�����;z�b����x#G��˧{�s��&��0��Q�%����+�	����sT�M�;��v�Q��d��<s��Q�v$Sص{6��t;��ǔ$U�p��s���;cFIR��{\n��H兛H�.�'�@)"{yepQ��؀lb��cnO=�^ޯ��zU���
Ѫ�nVv��Y6-�׆F-\����` 25�^>���uf{C�ߖ�r�n���I��"�d^�p2T�%	8!�R��Z�};Rw6V�r��G��z�﫚�Z/�RM��X_��8?H�
5Qi�U�ݻN���J�Љa��ª�vr1
A4`�Me�O?���=Ւu�)Vt�;a44������[j˃��2G�J��}����O:�k�x�?�h��
V��)>�WH_q��P�5��e�i�ɾ�P�����yT�bh>�W���lj9
�S8x��>�F��K2�O�=_�����y�L�&$�+���+��(֨�~y玎Q������.t���ǨkF)�쮊��x��b��l^BvB#ntGeTC�+,�z.Z����\I��h2���a`@o�cQ2U�e�C���v��K���׆?�jo-'2�S��X3��eNd�mԄ��������=̈́$�Y% �oUU#�_����H���n�h�oSy��p��ޢ�
a���.P��ɹÓ�'xYE�����-$�>��8@{��(}	c�,wPF^��{h4�� �,�,8k��yI� ��l2}1C� �s���4c��Qg1��W�
���|=���F�,l�Həq�!�I&.�@�ζ����dt�MREY�~����@"�r���"	@b�f������q�6�|C��2���Z���s����Վ�q��י���9��d>�(u��x4���I�Oe��|r%����&3�t���P��?5�M	YK�[	EZ�x�c[�~?��O<�K�M��\N���Q� ,D5�w���槑�G�Tq��L��ޢzl맷�������}����ǚ�݉"�(�0je+%��z������	>3yf��g�atT�;��݅	�L/@v�xá?��>޶�ɿw��g�<9�M�O7.��5�WC�ש�����l�N~%�5�}:�ٶ7Z�OS�#�h��;f��we��
���4G�:�4�H��
�8���T�㿫&A<�Vv���b���,[��Qq]И���7���n���	�/����[����v���Ω�J�,2��@�no�:,�UP=�I�9�w*4���B�{�5RЩ�)���b񙪁g0�p�-}wE͛�hwp@aZiU�fc	�Z�6u�*j��۸7A��#����m��EV㊋�U�'w�j����aN� IoM&��0�Z��C��d��\�V�8�ʃ�i��xa`~�!�џ�}�!M�K�%^� T��&�<�Dj�I:�B�7��&
҈G�(
�DaȢ�J��)�ë)hW%��H~#�f�7�^hC?�k���>:����O�@�Ts:G X�m�/JZ?���:��kI���n�g�w��l�I��!�y�C+#w�{��~�i�
�ݒ�u�
�gx�Y[�i�L�O? ��pJ��rHT}�~�:(��ƴ��һ��H��,>`��$��.�6�����ˌ�@5aBqnm7G�d��	��Ϟ.w%��?��E�;A1�n�p'�6��m��1�ft�^_	E��/rky;�[nPI�P�Kڎ�
�ǝ��}ŝ�c⾣.f��R�S��&��wa��r(ִ<�EnX�k��a�����y'����n���0]��mEo��>r����E��a�B�ѦW3��4��r�-�;oy��01�C	4��ܰp�V�nџݽ�mo�=m�ǃ��2~�.@�Xa�����8ɞ�M6UP��Jg� %���PPD�}Ba�l��m���I���e�%�&G�dk^S3�њ��\ 1�J��Z����;rTӑ���z��G����>]ke����֩
B'���8+O_��yu.�˲����+�%��B�Á�ھ�ܩ�Vc#D�o�h6 y�����>������s�Hx��n��^�c��+��{��/�$�k�]�Ҷ�9��M��`8k ��K�|��*��V��xC��W��9g1���C\��g��[�3�H��.<��0�\�&H3�'��ʆ[��lIg�Cq�����-آ��C��'6y��n#Sv���Λ��iܗ���n����=��Py�\�u���������+\�F�*63G���J�y|����Ф5��Ӕ���gH�?�O��
�r��Z���$J�p�*���3��4�E�RN�4Ǵ������s���+�Ep�M"��A�j�q��i��!��{�9o^��������iR�MlN;>��ޯWGw�*�SR&�y���r���W�*R۵�UO�+o�Et�_j��o6q	���+�K�a}�����@���_?��������#ӡ)��[��s�U�K�_�h��g3Å���c1�q$[BB�Z�Qm�'⯣�UDT>�[�+{Z�ax��0���^<����RRw@�7[�c|Xx���h�x�׳g���T-��Hd�}�P;���Rޖ�r:�~"|��(3�,8�M7�Қl��r�T# �0}a%��_+`R�ʪ�vR����H�M,F�(�y�[��2�;�X�K��xF���E���ӂp:*�E�N�u�f�wΟ�Z'ݙ���v��v�B7���*<Cp�~��(M>B�@��v`��9� �=�'�>�I�27D�#ZU� Jk��%����h	�K�g��2C-��DC!�������;8f�u �_gƗ�U�ҜuLܐ�7s���B�F�L�}֖��{ޜq�3��sRT:��-o]�@6BL>S���U�s�fvM� �����|b��1��G�`�r5g��
�s�5TAT���5@�&�@TNp�+Y�x���TM�&
Y^��p����~H���wn6��Km�T�p֔��qT	P^�̭�u��\�S����t	zl���%��:��g9�g�#�I�>,"�T�R�0�l���Qu�&��IW�튀��S�Os-��	w����oj�4+��v��c��Н03��Y"|�����QÑ�d&g�NK�*o���Õ������V�>�
����PO�ܬ~wi��H2���Z�x�vҤn�n�<�V��p�)_x?��N{��W�8�2��9�D��a��q�48�b@��N�B~�.��&���9 ��JJ,�Qؾ���[ q��:f�9{���H*�N���-%�J�8���D�txs�zV��UdJ���\�MStY9�M��V�<̆g@�I��� E�PD���H�ۉu~sb��u���H�L��8����U�3^�ּ� �Q�^E���-0�$�C��!�v{�=�!*�\���7I�c�<��`�|���q�M��e>�+l���b'Ʋ��*Ʈ�EO@n����]gҧ*�aw�p��z�������j/����+F[�w���.K�2_�m�s35��T�в��ʪ�xuG��+��Kǀ!���u��&ŷA�P�
;��~z���"����h�x��E�R�T���Y�vOL�4����$���`�Xu8�V�.���*&7o/KO=]�T��s���C�5Jv��4;�̈́�����]�����E��r�F\B�+�N?��&�O�r J�0�AܔG�";;�(����Fh8La9��������V�7����Ёti}��׻�>��ONщ��O���#|���X	!�F����<�.@n�>��y�~�I�%g|�_i���4�ː5����Gw�P;���Mȋ�?Ҕ9��v�Z+o�L�D��c����*g�o��db��ϠU�*]E�߯/(!gtXlt�揟�Y��b�׽���OC�Ļ�_�6�5RE?��ͻ����:��������)Ęy@��E�Qc��#�b��k��x�a�UN)�Ƽ��\G�u�~��a��T]��f��T:1�,�?��?��������};��{�� 0R�3�f��Ak��$����V��3�Iח84	����ɣ��`�`���%�MS�<t�����aA���x�YeRq��v��/��-u9�Q�,EJG���|���=��l<��ǚڅ�0̻�b�Hk�"���%ä��ʧ��zhgI+����ݪ�'{�͝�DW]l�W���f�i.ъyM/���/�z2���GZ����JF05�?��Ϙ�D���	�vu�N+q��P��m����>%\����(�,�WS���v�WAhV�B ����B�1.��D�K%KF~ƪ��Y\
��t�(�ߠa�d�{���<����_G�
���9����l���X����c��T��E]W�o��e=g-'�dc.uꪽÌ�!.Kr�it��O:G��6���Fߧ/�>���`�q;���/R�`pѠ_�B�I�!;?���l]�K$��dGf��1HO>PkE����1�%����֡��q?��m.���L"�Y"�G3ڙ*?�[K"Gx�z��8��8�R���Uʁ;y_��ni�(�.�㟒��Y`b^��P{'�s������C��5���&6nf���t�9���k�o��6��������[.�]s��p���>���='M���en�~�������]k��*M���MhH��q�Zͯ��a �֛^[�9T�f�h��}�%r���&�LY�-_��b� $v�}�A��L�6w/re�"���V=C0U�^��UȩiߍT~�6�'�Y�rr�ɾ��L�	�m�|Zl=b��y�)Q�h�%�W��SrQR���Ds�0x�v�+<�B��9b����T[=�E׀|:�eko|�CP�}vW, �%�SPy�#��P	��ѵ)��~TR����39-�*��Ű�C�J�ylv~tZ�']$͢Z�	r�5�I�s�q ́���«���	aմD���`�Q�,uN���&c��h>�r�������D�߉�ޮ�֦������p��N����z_[S!����
,
n�������YiF3�]jA~:\��U��-B���t�;��~i��Ϊ>٬�fi9�D���
�fv�|�U�Lc�-T�g�ڇ2r�%U��;3U-��$�%�F
��[�}3`��zĈ+���؝) ��	�]�f{G
�1��u������:�s��?E�ϟ�g�J���E�_�C�0�(9�H�[�%�Jz�TQX8c9�֚��8�I��4�1�H�;�<�Cx<+������~X��I�:��G�ʋ@k�s�Ƚ�U�W�5�j���H\�R�2�.��3�V� ��5��'�����2Ba �(��\����|��	�m�Ֆ�o[�qo��+�j����� n���bߖ��2�%w:�.A��9Yh��%*}+�_�>����!R��:7+T��|9.lև����D�C�Sd5�ĸ��<V_W"�m3�7��E�/��9�Y�����RiM٥����;�����6Ct ���,O�bD��]K�{�q��!�z�g�x��R ,KFt��}2��H�W�!�E~B̢�ݳ� Y��p�f�����o�ڧGA-�W�ڦyG�<����_7�ǒ�v��if�1�Ek}�:j���<�U �� ��Q�i(G�q����P�U!�P|Px`Ʈ��ch�E��WU�F= �a����	/�l� \K {rP���U�ݒ~�j<��Z�-"�t�9ɐkQUa�� 8ȱ�`�/b���QK��Z�Z�F�����I\��HE@e.�/�HsO��g�.��Q��:�J]�*�����ߚ���j�؏ۮ~Zk��}�V�@j{q����!3y"�D����31�vm��EO�o�8Y��3jcu8����D��2YX��m��b����?��'56v4��[|�L����6}5U���o���mLa6�U=�{Lk�B�j���Pu�D���w ηMsg�8�[�#�������C�d�0���#��?O����M�T|-A��I5��y�0�xY�Y�d0sA�&[*	��g�ʂ`�?��Z³�gD�?d�$�F4��Lg
�5~�)�[�W0�!e.q�[D��;<甎XV�����������[��:�e&�"���
1q�3a�����ݜ;�'t9���B�d��1�qȂ�	��G	ӽ����(��kq��9�s;!
��Ö+��<C�T�xGv�*�����dM��1T���̏�	;Bw��-Գs~��l���w���!��7o7U���<�߷!�cg=�l��en2������Y�ۙ�pu>�nRU�&Z��2�����ϵ�EhKC�&}�T;��3z�oil�ݡ��$�2����R]���ak�"瀄)�s�	ZQ���C;x���
t���ԯ��~�g��ev
H;�]��>7f�sK�7u� fdI͊(��GO8@�ڕXםMM�Ŝg.j����X��#ټa&RS��K�<�S&��MԱP�2�Ei�C������=�2��vf4�1�����p$���rJ�g\)e%��P�K�<�d6��O;�CK+&�3�sB���b�(+����w�K���Q>y�1i�y�T�ZBM�`���m���5�R繎�-^!oj�I������C�7�/9���c��
N����U ��:�����N�i/����Ek���Ӟ"�����:xL3���ܮ�������{jp��X~���˭G�hR�rjuF}h,����CЕy����U��Yk�n�Y �άʍ���1�ۙ���8Q�H4:;�oI� S�?�,�:�NE��]�`��q*���1
YP�v�f'-.�{@u�z��+�=67�YdJߖ��HY�%����F�`�IC��֖����ZG���f�Gg���n�إ�a:f�= )���DM^otLj�Kj3n_��&�x����	���'$��x�N݀3�/Nш�|�����c�o7f���X���T'}w�!�3�N[���;c�8���ˀ	ji�^���W�^�@�v�5���a����Ơ��I1���f�QɻM��E\��!�n��"-^�rgo����p*!|�a�obi'�!�G���+�7C�h���L+�&���<6n�"�C�а�����������?_T������������Cȅ.�hq��q0�-�1�x'��8����	�H�@��y��jz�_ZK�X�k�X���)\�"P�oI�!��j\�a�'�&�o	P��!�ĩ����!X����l��,h�WY��&�I��N�����U�?�����;Qe����8+��A&��^o����'��6���Ӥs�������0A�ËZA$�m�����u&�͙��/ϕ�7��/�t��l0��߈0��M�)��5q��J2f��an]�r�1�׍�èHJ /	os4L��J9E�2Y�^�n�m^�S	��.��Cߢ��7ʬ�F�J<�M���#m���	�e��K9q�N�s͊
�F��V��8_"��� r
�I��z���\g��5'@(<ՈQ2,�Ο;�4�8cl�J|���kK�D�p���۸�a��C�n��m0Ӌ��s��k�c��.
D�g������-���>��2? ,�Kg�����*�<�z�鹑+(E�-�;}�8C�Ҽ�0I�<Q��e��]GuX���ա�D�K��z� |�j��fBl!��ҭ8}��^�<HDP{�%��H3v���e���zNʅ~�Q#!G���t�ͱ�z��*1ROй�y�k�u�]�	����S���xc}D	Ո�&j������Rc�8�`���A�_�[5��a 83� ]�����;_V��=@너�uJ�e]j��2���M�hT^�0
����{с�Nv�1-Eo[�kV�"WC;��֤"��a#	�cJN�9�}�?*��m� �ZD��mY�Q0D�+i7~����g�v����㇘X���ǰ�(���!CJ$?�1Ǒ���}N��Q��y$�! ?x�~�_��u�	�����.4%�&���W�_���'���R���Ժ2��]l2q,f���hNp <{7��W�)����=�e�~'���x�B"?�(ё�M��iu���eU+��!%��LM�풗n��� �XxуX`�0�vF>�\D� T�|�
��K�*���Z�8uy�,���,;Bp��)��lթkPƐ�@H���D��h2�JūLҸ�m238ա�a�6��$�ժ&k��{N������c\�6@�4��Qge��F�;�ɿi�><��WW�s��8L����\A���3s6��l,6��ȷ�b@pǲI�QC)���D`sJ��
��1�M=Li;�T/}��4똖r)5qo��J�-Ƞ��뵀�~A����N��j=}>�	�k#f� 1��^HSaK���>о~����܌Op�hXvf���a��_hNX-�o2s������h�m�����_C��� Xp�����-6u�I�j��ץ�fu���=@џ4� {�}a4qclVJ�p։݊^�?$�Y#��� (���+u��Pǫ׷{៙�8����%�j���� �@͡Y�8A�g�0�;�0w��\R��$�[�<���o��������9��E��K��Я�R,ڭ���M��@�ݺ.aH�k>��D���!�|Zf�k2��#�Ԣ�qZ�C;23�
�]�)��������+�Ӌ-��F��!��d;bo1�qp;J.�ʙaW�DNy��[�N3Mۖ��lŪ@�.�/Ps�
7Y��@n��T��ie��/RP�f*f����G��u>�F��!�Wz�Q���X%�� =��C��E�G�K��	ڃ��M�yԹmu�J��tYO�d��rB~c���Iƃ�j��[�0�K+�t�w��Q.�o���e��ݟ;�4�^@�-;�D�V���	kc?+ !�l��'�/��G��hX�P���\�t�K.��T�U�9��PHp���vd��ġ�Nlܪ��]o@���g�DA��0>^x��
���m�����Q&9��I��1pA8&�i���落�6~4�|o,̗\�I�G6��";b�3w���y�:��Hս:I�W�����<	2@��nò�����n�Q�$���C
1��k�E�s5��Uyѱ�$,i��~���ɖ5��\/��gq$uź�����e�t��xn]F���,���.�J� �����PJ�-l�1���>}*G0FujRR	'a�6eh9���+y�[����ZG����(uW���q��q{/�� i�Z�SWb���<�w1Kú�/������:��Ѥn�0�"GN�,���(�-��3�<l,�S�|���(P�|,�-mBޓg����Na�3;LkK���2�}��?=]~<sW�1ahVf�4{o��ͷ�I�W/�]�����d�b��B��~��<�Э�����ߣ?Z�0��T��rY���)�F=r׹V"j��mƟ��d�e�XKU&���k߼/�b�N�p���cM�?��ύ�>���sr`e���~A!�Y4���3����O�?p�/�*{����כD))I�s��������r���ᛱ�
�qF�����gyR����<�B�E�p�x�����'�N673�8��ȉ֋:T�$�m��τhZ�<;�6�Ga�</f��B��?̅?։y-�Lp�ZX5�%ij*�������L٦qU�,q��艱�4�(: ����{�?�?4����̿t�������(@��U>m�V��ǚg��m�}w�4��"3�62H����F��8y�-L��_�1�`\�YH% ����~\%КYoO��Z����]༺cC��U��L�:̤�������.���@��/b�JgB(wΦ�%��=̞yMFy9������{��a��"�W޶u�A��?&jlbp҂���n��lD�:�|��Q��%H3�V��i~L���m�����*��JM���+u����Z���AI~+$�ܯ���D`M�I�ci	@�)	d�o��f�xy�1�g�[�]Y2;#P2�	�%�=�Gi6��WFI�5?��?wMN0��ӡiỏ+pշbn8a�ݥO]v�g\��~R'?��i᫫�0���T8ţĽZ��+	B�/y���b:VǟۓR����y������t��k����l���J�i�̸g����3rR.����D	'����'K��/8qL�� j���+�uMR�XD|�˕3&� �%�����l�I��IM��AT��f���5�\ʾ��,�\LYp����U���!Ѫ�<ܣ��͇1�}�����.��C��h��T\��nB�� �����5�1,4crvO��WG����RW����ݩ��	á~R̭V�5�^b�$%
�p,Spr"����>��5��c@�0�')��c���7E���5!Ԩ�L[㗝��Ӊ�	���0]g~�H�G�]3�+��\�Jf��U��\���\S_ �Zے�9�P��\�4#��g4�rǡt�aN�H9/�t� ��"��� 	����P����6^���F�o��&N�k}G5h@X�忡̧���C�� l�}`H���iv@����afJ�{kk��y��46Ls�?��]d,]���xI�f�;�бO�w�@:����Iqu�x�*L��`�{;�E�kZԼ]���3�U's�U���k��MM˖�cv�(
Z��[o"��m=�O9Q���7k�A+#�D���![����c���Q5Z����?�J}�����/fԺ�
�m a'�d��nF�������9�)߯�f�'+�"Ù��D}�ޥ  �)�_�`��e �_�U�����U�z�͇���������FH���>w��Gp&������d�_���-���|7�	[��!�؆
��Dk�vcj�V��y �����zD�lن`>�ѷYO�J��x���x*n@��'b^x9Cm]Te��U��J��i�<��ɬ��@��:�������{��T')���͂�|%8%[���i��~�:HAD�ƂG���@����垡��EBǯ��dx����ǢU����q:AEO�(+v�8md-S��1��!�7�����'(~Owm�B�q� E��/ǖ=����om40h�8��.i߻�G���|o�	3�j\�I觑�_il�Dn�������#�ڽޘ!w/�¹�5&�RiЍ�d��W�L6�N�V��|-	��3~u=݋���:H�J#X�%�b�D)��"$N�
ɁF`�!�^3�$ၪ9	�]�'�y����b���� 1���'^s|R}.{<�G�3���a���~- ����Ȁ�˥-�I�c_aW�l��Um�~
J�P�_68m���˜G���+�f@��WWW꒎n�o��/�f�x�;�����d����$���]c��������&��p�������0��|(�}��ӂ8�V�A����'��'����_���%����e�"�r�Ua}��
�(C�E�o������Ć���}&�-�w�wDKL��~���Y]�����"h8��:��!���ۀ^�'xi억$��I()U�zE���1��M����P�L�/�<5ij9Cp~����w	����֖����p����ۆA�uxɧʫ/7��_���''zj��!�z�G��ѼiF�t�;����xd�m�� k��?R��dߘj���F+������x4/�	�i0�b(a]�$ɬ�P:�7��8�O*l��f.Š�e!��W;�>��y�C��24���}ҽiꊑ7V*6�0v����2[�A+���ʶ�,o����t��	�3���L
v�d�'C�ю��;�(�������|i*R&�T0��܁�zs��x�Y�����|�I���,�Udu;f�ȍ�q�Ҍ��WKu �~)%9]<�$1Q�8b��?�<?�f���K�po� ^�[��q���M����,�Td!d�Ԃ��(��Y�Y���@V�W��=�x =x�����"/������1�������
? � p#c6�ZUǪG9�\j����A'��xA��M+��Q|�?����p���e�7[bI��+�8o�(M�U��0?@5d��%&�/+�)��G�m[�G&V����FS��^����֬AAp{B�y���y�Y���q� w�DE�kF}��}Yz�Xc�t>^`�.y�Fc��S�/�AK��H���d��������5/�"�v$ux6�%�UO�xW��BƸ⥹=o���p�\��T'vT�8���]a�ʨ�9��4a�ط��k�O��T�k������Y(_|/H4���pJe�+�0�2��xngE���w�|Rt�<�f��'Y!�C�h@0�B�[�,�Zf^5�&�hx�6�/������������ꮅ2�,N���ђ���p���;�R]��o�M�����2\Jk��V77�d�zn�,�y��H�t�k�qo{�f�rޗ�<4����5**�W�a�p���Z(�˜�V��)�8����2h7=���V��&�H�QO������LUeߔ#d����Hr�?HZ�@�Ѡ���Z�	F>�t�$PmX�����e����շ[#,�@)*���	��/Yi���<k6��v�sz�(Y&��$��0M�jg�H���A$�����n��A�%nسVE��M����ݏ)���Y�k
� �aur��1���_;kzP��i��|w2��UM[��+���k�Ԡt�.����j9�|�$�M�_��76V��Py��@Ď�'��c3�n4tO(�(̍.���l�j�� j�g�xޝ�?��ؤ���k��ȹ�O��G3>ʋ�ԛE�	����Izg��84�������<.~���h]C�1��4�^���ƒ-�<Q�^0��=�S���CW�H�Ճ�vX�<����A�Z���zqڻR��59R[�����\�B�' |��7 hD�0�:��+��2�z~��1�o��a��A�>m���6�*�zE��)��(�&��r��|2f��{�;�axu�����������#�3=����m��#�N����u=��i��n�ՎB�����N�M�� ޹������i5(��1�4�z��w�U7|5Ԙ})�/#�v�Y�U�TK������>A:1P�2n&E!�}]p3�G���񧋿|o�M@������������
�Ӹ����1$l���N&�f/�w�T��=?gⰹ��*=(�5�������_��<�]H/0���s#�rD�=Y������M�Qh���:����?��@l���a�)���H��O���9�`ͥ�t1JV�s�`�y���JD|tѤ�����M�aff`�'�&�~w�v
��sT�O�6p+%�f��y*0�f���\8)IN�)�(Kݬ���@gF@����U�1��V�	�^�����Q�Ӝj�$�}�9jY�;f�1��T�Ua�~��9�C���Gl�P�f�]+�r�q������ ���Z���=)����"�7�@$���t�:gz�th�ԇ��&| ���H���i 3��x��p���iT�hH�_��M��A�o �#�*"=���vD�g��q5�#9�p�J����a��?J^=S �>P��C��� H�Ձi��&�f���{S�%+���F�����"lvܳP���TD����q��gyZoO�¯p1����W��yhz��M'AK��Dx�Q�iU����N>�
�	���cJJ,A����ưJs���v�����Ű�¼���'J�nPg��}�H꽷��Y(򍿄16�;t'���p���W��Я%U�+U��3q��sO����|2'F��f47�*Ie�o=���02D���3��\{6;K�i�u�iU�'��ߍ�*!REP�$�Ee�Jb_��Q/���r���|)4����k��7��q��l�QW4z�1���u��v�:��3R�AX�RC_Y||DU}�Os�����!5�RTy��b*�.nP��k�2ғp�_6_����ߔM�Z�c�Y��y�Dk��Z��ZV�����]�[5�g�K��#�^�e׊�ƞ���z)�2eOg�E�8��;均�����͵d��������Ceqm�'g��@�X��}e �T�0T��-?����,݄GT8 Ts4V��?q͗d�Q�NQr�Pw�sW-�xr}$>�}v*��y2��5V}�ߝU붺)"���U��(�ng�� �����\e��a.xD^��ho�T�y}+�.���%��qK��Ej����d�E����̃�:�o4�Ev<2ҏ+��M���Ku1)�/���4Q}�Ƒ�0�l$����_"a�;" iq !`A�<f�{����=��r���~��"'Ja�g�{�p�s��' �����
HϺ. �ZyqZ�|�"��Vi�0��,:ΎF�����p3jF��޷�Po.('��:"$�{�[�x����@4SM_�(�?�����R����_�����BM�8<�f[_[x��k��.��[��-���B3"N�.�;pL�#��<����R��x)!Ķe\�A{��J9���M�c`9<�f�g����徭`��yz�VpB�u���m�8�zס9���,���W{�j
�Y�
���rl��?�TT�� ÃU�jP��.kM;�yd��z���շ�i��S��,�J�=>�#���<��Ͼ#ѯ����p�䜠̯��wI��0�ldN�f�ҡ��d�ڑ\>B��|�ɢ�u�_��ʝ�"��^�u�h {�g#�E*�u������/����m�6i���k�#d<T!��y%97��'Ɣ)��w���e�hC���Np���U10���T�3����*磺{����JPF	�����v^i�;��.op��i�[?���!�$�A�����ky�����!�P����L���V���'�g �B��k](���'���ppvwǷݑE����1�et�S)���׭�C	�o��B՗bk�O��8�M���R��ڨ�a�����R�\cp���U(Ѷ,�I��a�B����$�;^����e~]v��h�D�hˊl����%���8l ����0M������h��x�<���N�E���^�
����;������(/Z�Y�����vhrM�زcV�Z@�R/0���\x�1�+ޠ.�mn�XxE���y��>�?F7U�����~^�� m�r.��m������[׮E!�s�re ��)Y�ӣ[(=�@�$8��H�=�9�aSMR�*'�T�QZ�fE����
^ g��ؕ���	��U�ƒ�
��K��Wz.�H��?��
��3��J�!�i̶`����x�}���A��+n����s�K�t��'�����%[)�L,B���U-����4 t�F�_��?���������e8�$
p��7�ĝp���\l�a�1�h�좰�}�E@��?���D:&�nZ�n �o����)d���X�X�"�e��ʍ�e����m@[zL�;�y�~_��Vc�;�mY�(�LM�#�'�� �'��s���9����q����t�b%�Yn����1�ݰ2�.����5xK�\ʮVY��U?��i��s�Ǧ ���=����;|�hPJ3k����Q1���������jE$׃�
����.,��5��;;�&̓�Ѳ�$_��=ǵӎ�\cQ�yP`Q6������܀.3�lԳ�\%j�Bz��*��[�J��MTʵ�g�%7�j=�&�=�ņ�m.���E)����1P4��8#�Ŭ���e�@k*�φ��P�4���Jøp�q�aA�Ѫ�!z�|Jjz�G|�P*����;���a�-1��eY[m;H�+pn�
��n߈�uU�\& ��jU�k�D�WM���QS�Ƌ�rm�vu�тOc8�����^:��F��NϏt�����*�cKs)� B_$o�W�x]��!3�B�8?��##dJ6!EK��ȩ^�Z���:��t]b���Z�ƪ��t��8�J���KP�(b����)�H/�_yA;�w�=�א�f�:�s\P�Z��q��sԀ�u���f��L����뮹r�v�/q|3L����£|���&�#�L��|:�HZUxz�AH��$K�O�{A�0$T����#�,���&y���Q7��<jZ<�H�J��%�}��i���D'H-,5�Q�X;,�����@�<Y�����.rs�:l��Х��3b�-`���+�%C7i�3���&��T��eaZ��6!�ZxkF�����|�^5}�S�Q�:�-Z�p�9*���y��.1S!��;=���2mZ#v��c�,�V�XmF���h��!8*~,#�13�{�(ŶF���i��G`�o�n'K9�H@R���)�� *\�+b��v��\=����_� t������/�s���X}����-�Ip���&�@��y��K8K��YQi�b�k'��*NT���j�9���V�ķ��ܤԓ/�U����7״Y�l�r��k���sjٹ�<��+f� � [�����.�C���Urĩ�����e�������yϱ?3�ߐ�T?e����C9� Pw:�D�B�]���O��t/(��n2�?5�{��3��rT�s�c2I����h@�������H�-v:/[��h,�UIe�Y�@��kų�.��
�[�:��KOU�,0�T�T��L������V�,��n�qT?x��bl��-��
V�j��O1��͸z�C�܂�Bc��2�S�E2!�T#ڎ��r��39��es�|=d�5о��-enL ��~P�\&�Yo#�v� �P�Sz; �-*�ƛ%��k���Q�;��S�"�?a���w�"(�Ҭb�'��
�{X|�N�}W����O���J���̴/1c��Nq��0�h�}���c��$S҅�Q^����te���S_JaFl��T2�����[��Qm �gF��E�� +�d<c��u�x��Q��z9.W�"�)t�P����!��~1��!���m�)@S���=&5�˼]KQ�?Koҷ+�л�F��>���1��6�m��%E=�/[h�	��q�ЇŃ΀��eJ��rC���.�r�,�U�8q��LB*�V�_&��@P���6r����T:B�+i+[C�CCGm��҈�kw��T�H��J&t\��r�do�;7�M�Bط�2�{�$����h����X5>��}�.��1͂�(Nl!l��v�r�O��Ȓ�i��"+`��{ jm2B�DN03��\s7�����>��Ac�;g���)N'������p���ӟ�4������ro��i����ٚ�T�J�<�$J�T�?�7;���s�9p��|ڣ��ɨ�)5D5:�ҒȷC`�M}���-�7"�".�B�/��&ǓF�>:�j*�:TL��]hj/��M���:9�D7G��N,����X���+c��vi9f�;�����p�$fH#�ȳ���ހX/�=W��K����tK6F �(�[DJ�-�Fc��7"��y$��\����)Nd�r��Z	�G�vv� U��
y��~�H�g�ȬG��w�ʊg��<������!|�C(u����^�^ڐk��b��t�!�G�x�L�϶���Q���]C�*O�d�"ȇH5"d\r��NvH� .C-��Ht� �SXI|Sa�_#Q.y���7�!ʋ�%L�it�$K,,��U�%o8�|`9�njN�sC˿
~H��G������,���=��+���ś��E�J��դ�����.�#B�Ӄ0i���Y?wnXR��O����~�lfQ���w9���'�sϩ{��H6�c���c����qE��)���B��F��^��G�E%�u.0+�r�6"�B5&���|qƦ��HU���5����IٜN��)J�8)6
��o�o��R]�e�� r�X�M�̋����|ܥ�AĠ(}��d���PE?��pQ#�OG�&���S��x�����(0f�g�fq�����>�=Zl$�6��d��2^-��oJ���p�8;0�;��� ^��:z���spC0*�^�&�i���U�/
�7��z�,����^��Bu���W�^J����)q*�s�������U�蝶I��cDpXq��|���a+%]�x��$)[^�}���=C��y�z#i�`�l�4i��'�v��׼˭r�����#�)�s@��Z�{2}�6�L�i�Z����w㢞��#���,�����ǟ������#,�Aɵ83=&Vʷl�G�E)������f�w��؉���.l�@!Ԥb���نϢ��
Mc���묝�����/hņmތ}iϙ�9�7��Q_�x��/x7�.+�k�ڀ������C|���J��y�x����.[9维��O��.��,�)"C�͋(�#,��������(A�w�J1f-�6RW�Yݬ���V���1~��7]lx%_�IvH���������c�c�%���C[K�I�w�J��&0����V?4�G���/8�ު��ҎN�0�����R��qQ3�a���z�rU!��]P�bp<���S<�pV��t��LA�0���L��_nU�"э�^zU�GM�C�\���� 2\��%I�İ�'�̓��)����N����ݟ��ˠ�0�����x"uB}���h�SR�T�~� �r9�ⷄ��]�@TP��qsc�`k*d� �Ҏ	�",[�VS��X�3m�K2�&�u'c6Uy��h���r�C��#�8�֜'~K�e�H�%�!�Z%��g�J�blY4x�%+�O�{;$cܨB�u= j]�(-��ې-T)��o�����p�t�׊J�
ݩ��FF��z�ԃ�2����23��m��c
�]7(��H��2�^��ZK�.����/i��L��(ak��/�FS��W��pB�W�\p����, =��3�Ln藧���w���s��  ���3���ݞ
���˨������� �\����@#ּ��LrZ
JR��.�_���֢!�h"O���N���~�b8��u�=>M��\*N �G��!4������P�,~.��wa�Ytli�� ���25`��?�}.j�r�K�w��r�v�+�N�	7���&�ۨ�b�5��<+�o.'���&�c��!�r�1��e/�;���S@hyՅ���R���Ʊ��]D⊕s�8��XS�Њ?g>�$�.1�Q���A���{�s�0�Z4C�߫�5#D2��o!��9ڎ�ٶ6mxՏ��⪎�a,NJM��u�.)[����s
�:W���dEYO9���7ݥ?G|(��u��	��A̍��r���;��4����z�T�*��� <*P�n�!
�0�����p=�K���iدpx/������򗁋��2�����0T���~�B����C�����sӽ���R�:�U��-�;����B)x"�#HU᭜��yƋ�����ɽy�����h���Ca�1;�V8ZZ��z�5�oED�	�T�QG��a� B�S�0���Uc��Z��rT�SA����NB�Xr��*q��.�YP����D|U0�c�n'�q���Fj:��+c�
l䯵���l��e.�V�a-_X߳��y'�6��&Ȳ��b�օL���p)�gW.�
�oP�ê�g0�}LȈ 6�GFѴd(���b�j��$;9劍��T�
&G�}L"CH��F���;^��&B�&�2���i��=츌�(��}�� �|w$v`r<�-��Ky��w��AR��܉u���5��x:vzsh"݄x)��.K�~�R�瞎 eu��o�Y������d=:}4�|gJ�!YW)� e�>
�OO��]���x|yO؇sQ��]�����a�Gk�I�[E�6�~� �w�U�u 3�������T�s,�ۼ�wa�7��5.���Xξ��A��|�G�Q߳����g[6F�B�m8�z�j��y雿Q�rN�M\@�6o�Q�g��1�#^[�+���DYd�!�1�����I�Z{k�z=��u��E�>!MR�y��w'6��v���8��' tR�O�0v�;�OE},(/!~
����qФ2jƤ�>r���[+�����l0�D���q3<D%�B�\�QK���&±D}1~�!?��s��L{�;P%S�+ݥ�vv�I�m���a��:#���)�6"LK�4],�V9�2��/�(s������G�+1�+Hm��LL��3�N)����?<O�Yn��3�$S�I��t*�>��ܪ�j����H�K�\kk{�r]�7UΆ|e���_}+(��OyO�T�)�Z�f�J��Hq<�U��xۮ�w|E�y;U.:��G��Yo�>~q^'���k4��S�y7;���U��q�sT��n�ـnQ�<��`#2)��^�F�� ��ۯ�ku�
�/T���H~��PVTC 8��$f��/v�2�4���S��r:���y�LmkƲ.y�u.�gU��M�6��M������4d�53mw-T�ڮ,*��Fy���y��6�^;��G\=��`��!���hRm�Rl9��]'8w���LH֛,�8"W����ݨR�����Ș[�9�z��,q��"R���@�x�Q���%w+�g��Ў��pVd�V�Yt�[(��:�c�B�i�-��\����!��Ѭ�R��O	�gCua����A����¿K�Fi.�O��[���7��w>_����j�a?~ �p��q���`[��n��a��RK7�ěQb�ټ\���~�G
���������ٕ���@lxUjQ�[��TeD��z 隿l/��5c:�����,+�dI��uM/��)-��z��h���Kb�8a��7��aC./��I��klDJ�gz�5���g��zu�,���YQ%D#,�v��L�+*���_�a��"#E��h0J]g�f�$�����W2,��J����(Bc@�"`�y�^�����g�5�����E]y�+�����!�5�M�̅�Ψ0tâz�Dݙ���_O�(�ᢦx1+�Mo�ܨkX��ςI��#���pd��e4qL�>?�Ug��z����n���G��aeKqP�a�72D�Z�e�<_g_7!һw���g3�/�iB��ĕ�k��0O]�0r��s�����0r��A���#�H��3�$/�JD�d�\a	T���xw�[H��o~Qw�7vFVch���wԔ�nɔA�9��d0\3�5
v�5n'V/-mD$aԽ�C��θ;�}�x@����uz�9��N��X�������Y8p�q�Yu��l��|1=U���A��k@ �2D�s��Hn��hm��K<}W�ڣ��7���;����Tz\]|&6H�àn��m��PK,ǡ�ӭr�G�,��7�,��R6��������וn��`z����ь8U<&;YYe��c�3y��	��Ne�VO
�7}%�c�Ki�Z����<zԎm���]<��+vc�v�Mj󲑆�li�B�JW�{���g��0�9��{`;�'�""7��������;�Xn��f*h��N��n%�/��8Fɇu+�ޢ1�P�RWͅ�@_)9�\u�m?5�Lӆ*��@v�Jj�)R��d����`��hrAˀ9����c��T�;�5�VS�%=S�"@:����`�M����Tz��?�,w�S�w��cmG=>"�q�F�ua5�U�#]���c
�!�>�cC�lڻ�ED|:N�vP��SG%��Y���X���#�N��C�v�#
�A�9��MJt�)��G&�'����Y`|��2��y4@qS)p��:X�۫�.����P��izd|I\x^�*��y�ҟ�֘֒9yP�=i�(�&{���G�����_��B��x���/��eX_��S49��i>��}X7�yjYZ8^�WRL�E,��9��?嶿G�����]T+ũ%Mu͔iy��sٴ��%������_�UQ�W�6΁=���ٵ	S�Z�g�ԓ~ ۠�m�Fo5b�	/���RN�h�c�G�H0Ē�H�MΒu�q�i9��($��"��4��ٯ�P�sx��<�\ζ�c�y�peJ	i��k*�*I6��o���Ң����q�N�0D-��|A�\�� `a��n����	]9FG"���}�)��+�[A�%��b��3�g��w^�Њ���g�#����L��s^�ː��oX�1��5�s�ۄ�:qn[��.#wɣ� r�^bp����f@�w�ee/�v6����Y{�]�qH1��û;)+ 1}�����Çh�cLʚ��dؤg�H�_m���'�꫖�S�~���q*\?��b��!2^��L#�F�#�\K�����ݲ�f�Z=��r���[�����g�?��}���iɘ�ň������e߄��1�O�o�q ����8�J��-���&��%A�R�U���n��:LX�g�.j��݋�����^��w��w��= iY�Ag0q�ܗ��s$k���R�̾!}G�@�l�
:K<�\��U�����b�mM𨊔�U?J^���V�;��e<�@�{�
6\0�4H�ྦ&ܗ��k���C�����ĩvb���9�Pd����(�=SX-�x7h�5$J�!��?o�æ�Q��a��� O��O��
Pj�w��B&O��a~��,�H��τ�� %�d��tRb{��!�T�L�s�3��hjW�%HǌDd,�m��6H#y��x�c,����W{ �z��˖fm����A�@9?#%���=#�
��접�j2@W�OS��3N�"d��ÒicF�����i�v�"�)������9��5��y����e������fG.fJ�z�+}1��M���^�I�.|�;��]E��3)��R��,G	��+�ړ�:�y���| �y�\�3�|��V��@�҂��j�mwJ
�
��5�a0�JG%π��M:��Qؘ~����ޢ(?s��85�� ����O	�Q�eCANt��m�_z/&�/ﶸd�7\Q�45�x���I�X���<[�����\U���;4�@#hKR�LV,��k&<�NKd5�3���������l[q��R:R�����z8�����Yp�@�݂^�+U*���C������>��B۔S�ڭ���[}m���gY�/������3�N�HI���C�t`J*��lk:%Ɍc�|����'˱w;�i�	��^�*aR�y����Etd��!��f�e]l}*���R��	��m�n˘�|a!�1�p=|b7��lx�?��]g]<����V'���u�ϦXK�l��Is��m=���P��`'"%?�n��~�b�����1T�X�Η\�h��r�_���C_���wUc��ޛ��NK��f��5f�E�5�g��4�0R-ʝOJ:��c��=���l���M�v�8�hA�^y>��+��o� <���u"jy�8�W��@�ɜw,ۑo�P� �מe��a��XU��毻��;R~�� 9B���`e7�G��f���M�2z�,���!N���I�����R*Ha_&W�!�X^}vv��'ڣ�10y�v̈J ����l��o,��}��xT���0�/���2��I�nq-���g���,yJ(9��Z���љ���0j�I9�0����s��}! ��ᗛ�̃*���v�O5ˈ���k��5�fn���uE�Ah
%��Ҹ�	���s�ڞO>�w� �@�}E�������C����A� xT�pϓx���D�ߦ��+�"��������w5�/�ƪ�������M��һV��q����
U3�6�i%(�G��挟�u*_:-����oC�m+��	m���e�����m '�<� ���>).m!�_�^���\)W�`�A-����ڞ��\j�>�c�qmF�C)��Ʀ��w�l�V,�$�&��(��D[��ߡ���g���s�s��F8#�*9+Q~�J�S�{P�nk:!@U����~cZ�:�l��j��0d��6UR���Ye���p�K��΂`I�~�v|��l�ۗ�к���������*'S�}2��b$����d����rݴK�=;����bR̙�.
�vCJ��c���͛��� X���]���2Zi�]���[2��ʍ
�@A@2� ��3�C]Pу��?yk�ݐ`�fvP�X`ʺ�	��1�x�W��
��PtzO� ���4,ޗPdp��)��#H���3l�킮���t��U�3c��_�WL*&Rˊ8p�޿���hU*Y�����9��?�МFߵ�;��2�����VyT�C�%���a(������V���Ջ�枿\i,��B�sF��nS�.�3��mC�B��3�M�ET��1U��}`.,�頖��]�(_o9�M}�e�
S�����{?� �ğZ�,^�t'
�r��e�_����r��(�SВ6��!6�~�Oa���*2in�:߆,5B�شN��cA�]+v��P��R�vH��
��n����Y1�d�r-hē>9��fv�����IkO��NY��H�S�T2F���!�B�^�@6�:�\
*�����;�rb5˴S��C_���m����u��R�� >-��aG����
ys�I4Jv8|Z",�Y%�U,���ƪ�2�M� �%^4��w��Ϯ��Ȯ�t/htai�}S�@N�t�6
5B��m�(?{��,Smo�{�7�cl����ݝR�s�Q|ya�;�V"��ꒀv��S�<ve���ؽʴz���fRaw�T5��h���*�|ǈ6=��&8��ړ璜v�V�SD�O���6 n�A�6�ʚU���C�H��C�Fq���#�OZ®]vbx� .��Nt���M�r�L���u]_��Q�C���[b��
�����&�uܪ�c�S�s�[H�͟���wBLg@�AP꣏r�ʿbw�4�$�>Y�	|Jcs��S��s{�l&>��+c-�*�w��D;@��9��I�!�4 ʟ���nn
e�1�U~9�f�;� ��oNu�;��$Hl��/�:8ĩӟ�ꔂ�u��Y��I��z���c�oWm�<vt��M�q�2QǲuU���uS��ku�9C�Z�*O�����|�k8�����]�C���o��<���#�'�}(�.�F�	Yak��>Xz���������;T�I��\[�E��0{�qRG;F�m]��Z�%�g�+x��꟪�7����n A����K�q`W� �{����+Q/��s�[ѵX����M��Sɔ+A���Z��TCc�L�?|i��w/;�7��$}3���A\=�����ג��K����2F�g��$c��.�x��Zd!��U`>��>@2M�"�|���9�0�.dH }�R:t� 
��j�8����j[n}ZkH�����!�"t�)p솨�	���qh�T�7�ք�.&�^�ek����(�V��a���()���EC��ݵWO�YM�cI���~/��a�qZ���ޘ Hq�EЪ�	�uݜ|���l�W��tɁ�1|a7J����5��
��+$c�W[�g�4��5\�p�T��YG}�K�GUA�ߙ��cy�TQ
�=�*!n�&cE�R��alA�3M!��&��s%;D� �b#��s%���S'{=�h
uz�?�S�U��.<��S��|��f��5��<ۑ:!��}������S��Q@
��u�8��]������:�1��H��C�@4�u��h4���BT^�Њe_r�q!W.�g*��1TV�FZ
�gƑO�S��q>���V`���ò%��8U������]ر]S�Cg�m���})�bxn!��$lW_UN�WP�q5[0r_?�R� ��m�ۦĂN&e;�O�d|�&j �W���X�Wr��S4�x��?�D1Ky����c�FV0^wĝD�<(;��M�v��HY3#�1u&~��7+]���*���IᶯQ�PY�֟�;z(u9k����"Q�y���􃨪;hX߻<{
օ��O��7r�˅�������J���KTOd��[��p���I�z�ęq��{v�*�?ҥ��ܜR���M-�݃���3j'�:1��X�%~+�O ��]|�7& ��$�Y!%��#T٧	�F������C7�6�\��SoC��A���`e�t_��٬VBk9c��2���A�B���[�]ڙ���W��^�����8��w\<�ɑO���|$���W�U]<�./��-K�o8��r��Y�Z�^'��&
:�>4�ʇ�,�4
��@�ɥ"��J����zm)3H�7��Ic�O�Z��q(� �Y:��n�D/;�,����N����g��Y�}���s9��"���c<!�+�HNJ���h^�Z�#o���y��\�����!�埚@�0��R�D��X#!�F׊��{'3�5��g\1|򒙴VJ,�{����8�axW,�4ta߳�UH��F�S��{�C$w�����)�/��.��5���c�j�4��ꄶ�a����%i࿹b�}�g�s�������HaCe̮_�X���3c����{>9�!�]w���5^��nj�eZK���W�c�I6�]�s˨ �hw�+]���LI����d~ۿ��8�DRE�xg��z�������moQ,� &��*��Bs?�`��<~H�;����h���X� ��F�!C?9���h��Q�PbE	b�4�c��}AY����䯀?�"��mٸ<�$7_�2��i�Bv�f�\t�.~h�]`��n�z�{{����l����.Nvpa���U**�����ˊ�@��L�,6�rR����.�ı�<�J"�^--�I�^�&�
=\OӇ�i�����f<$0u�nѿ���6��V�|�b�Z����*��'��I�M�ynz
��4W�N`�!�3��|h;+���d�$���a�俌T�c�PP��;�Ai� iF�|��l���"����EO��%0m&qsc����2
��#�$�K�������E�.6gZ?�8�08_�ԈȾ�8�Ä=�&�%)�m��}��X'����~�Vv|��}z&�=��0s�����6����	 �0=9��-jň+2j/)�ed4���9����ɩjW^I�������y�|�?���������&N�/��!� +6`��Y/+ڶt���)'��J+M�0Ԇa�n^����\�X=���J�j��/NS}.o�ѕ;02ׁ܆�e0FW􏒳�Ӂ[����� A=��E������1Q��W�������4g��J��4G�����5�c� �RM��{�V)���������e"c��W�+��h7uI�� �M���<_T�����d�Z��/,���H�v4I_���PQ�k?Ov��a�5��d$��"�AsP�R��p.�^�����J� ����S��T���)k�eߺ�:�B0�w�:�x<K -�őv�#����>p_b�A���0{��'�Y�H±	RΠ��#_�,9d����9 ��/�j�[T����xiT�����,!Z1��#�h4=�YMe=�ӈ��LW#w
��t��_��-(+.��5�}��T����y�:��H�-u�?�����5��`S6����-���v��\��sp噟۸�
���^�6�G�� �����X��@�[Ԕ���xJ���Ջ^x�7c�o�
��,�_^BD�����Ç�d=?�D0≭X{��O�����mW���o]�Rh��f�z�`��޸X�2O��oy�I5�)u��I�;�X8�(jUvt��� ]���D���rD�0	r	K�������~�b7ӓ����.�r���aޫH��_;MB��]�>�����sb�Z�5iHնh&��1K��?�VE�$b_�5u�J��zAQ�L��Ez�/W"De;��z��D@KX��|!�FD�k��<��a8t�o���=�l�mf�­���!3�|�ϊ
6z�]�c��D@9��&��#*��U; $)9��`[m��lE�'�` fX�)�w���`��)��RV�B;Eϊ�J�!t1.�Ƴ�pL����V�y�J����$YV�e8���	)x��Z\�@/o��@=n ��wm�8�e[)	��v�EȖ{YKh�i�#��8����^�AQ��0��ƦX�P��c�d�皧�+�M���S!=z�#�H�HR��#��Z>��#���@dxS���p�z؁�śU���9�g�1E��A<�z/}�A�L���C�z��f��hF4��
AXݕv�巍E��aW�<��
3/cQrU���Ζ�Ё�e˗J\� ����s��Z�Dz�͗��n��#�!o9K�G؄2��Y���[A1�2Y�-EV+KʧÀ�3wܻ�O�.��ZB+7�`_��\b�4$�����am��=:�����(�H`�.�V��'92���&;�]ķ㶫yZD`c�v }ֳeSX�k	����ueB�)rc�^��qd�-)�ك=v�dY.1�n�u���xU�Ḁ�] 
x/Q�鷡����AKn)5��cWK�	�L/䜋&�E�l�V��6�n��rSE�P&8l��*���p/)��9���?˾.��� f�m���-��\���;�E}�&r ��֦�dp�"y�v���/Sz+}����>�c���qıs(��$𗄅v@�>��	R�I��1�wn=�@?�g�V3	��P'I1
�k��@V:��,#����R��AC#V�3�<Dx�-��|�s��!6vYǝ��04�}���\��m8�j�g#�
UXxC��J*�h�)Z���=|��o[��o�����gԲ�b�L,�Y LA����u����:c4���ro\<*$d����L�u�|�@#ù����n��|�u�*�w�nLU�d0�.L �m����@;�P��Ok]�C���c��l4>�晞bf��}����z��eP��k���ӓmQT�o!X�[ę�Q%�O.��� 
��r?�:�a���Ɔ�-�R�.!�P}�8z���]�#^Y5N淠ݖ?->�Co��y<,��8�^(��o6M�qC��>��ַ@�
��H��L����O��*mXpw�ɞS�l%�G/������B^4�D�K��OVʕ_��!l3j�sǍ��e��~|$��7��T������$Щ��%H�J��������r��͊��
	��6�(ԗ�s|P}���f�"���ch����ьk�y�P˼��Λ�i �-�b�VxqO�F��N�Yh@QO���uW??�A
��F4>4��y�3e���?�$#|p�#m����k@bM'���ґ �Z!M3������B�/a6�'�R�e�� �Z�'� h�jkYZP&�5�=�hV��P�[��׆l�T#�h�'�>D��
x�6���M}侴���[���L2�{�WZ~!�:@�ɠ/r�f�L�Prܛ����Q����8leU�Z=��>�HXt�A7��ġ[�x���{�ut�"� ��b����ܖ�
7�g�=�L-�U��*ŀ4;~�/yP�H�Mƞ�UVN�s�(��G�
�xu�?�����'.��������~K�A���OEP�-S��NA֑�|]bl��a�q�H>����.j��/�M��'�~������!�<\�'�0��f+6/^>L������Y��Ɣ?����*�e� �����t�䇿i���v"���փu�N�'V��S�,�PB�{"d��r��C��]$��y�@w�j�*����e��;6X&TRd�����{�{���f��eA��%�EH���+ѯ揹�`L�`��
�)W��R�vC1账�^.G,� G`��`Ѻ��]' t%��1���"w�֯��C�l;;�i��,��iI'�M���1�=�kT�.Qd�/P��
��W2��(^���n\( ������R�����ETCĎQ�z�� ��:,�ŒŹz�Z��t� P�_|�q�4���җ�뭧+kn�l���]�OW�?�Qt^�"�䙈.o�־�䬲R4}}��!�H��6�
�%ˋ��E[W�!h�ˬ�s���e[�>�m����=�l..{a��=p��g��'J��˃�M�s��<;w
��bK���R�;h��e� �Z;��o������۴��y5�_�nF�C%Z�&�B%"���]��d�ʺ�X�r,��zg�t�';������ ���w
�C�#B�6NIƿu��U;%Ѻ�ē��r�zB����Fok��xp�y8�f�f���
]��oѠ��ic���*�	�&��P��>6�D:r�@��ʸ��^p܃_1@�JU2�U�ŭ�b��Z#����aa�M�:���+�삺S	���W�/�$
0d�9|���㵞��f�h����ΰTX_̾���SH���NQt�P�:TD�֭�r���&te�?WG��h�������ebRgT,cd�� 2b8k~`�p���"͈Do��C�6�zs"-�#D�*&���d}�d�s�e�/�ی���n��o2����<��aATF�yGT�wr���W�r��p��y�b�[U�cr�>؄��0�gY��4#���J�3�I�w���	V󈙄��=.����#��S�6�(�$���\ة]�e��Ĺ=����<z�	"?8u���Z�b3YS�(�5��j���	�: ��	�� m�s�+���ktlַl<q�6��$Op0�e�r"҅öt+��8/-i���S#@J������+"�����~�������K����m���T���8"���(�S���8(lZ�5��l%�SЦ��������;mȅrF�:����bje��>���8�)�ޤO!�~������nxk5Ξ�e�+��L���2c��M�q����Clw��p��A��]ƷL)�*���Q��w4�
e�ϟ%w�@�Y�/KM�"m5���������en�/�n�\�o�3��k�r�� Ж=t��ǖ�k�~��}�~�H4��^�	���䳨xÇ�Jͼ� �4��"kg�������ȕ[(IBP�����Ņ�]̔8iߍ}7�n#�Y���\�qӝ)߄r ��Q����NQ圾,dT��Ů1�HFlǤ���!��:����$�YJ��o˟�AK������Ɂ*b^"�@���:]�� �f�Rn���2�Ƈ
1c���^ݳ<z��DE�7�_��Q��\/���L�NSq�GĬ�^sT�����B���ZNC^� ��&�fn�����$�S�,�4>;Rr(��﷿��PJn2��>����t���P2�avȝ�q��߽/�<X�̎_&b�c�� �N��q�b�s���Pjĭ���G>«����7��8��%!�_7��A�sD�?I�:���.z�2.��x�ʕr�� ���W��*�m?��靑3����̹�T�^���&h�(Ԉ�r����b(��(��^u/>8��x}�Y��phXa�"�q�l���x���; :]��>��-���f����6�̩l����Aq�ڞ�	j"��!�f�;*o�_�h�x��* @3�3�*"�* x�3㦚�5���K��9�06g������ْ���[�u-��{M����W���c��v�;����^�8�8���g]mߒp3�Z$&�U6'vo�Q�#k�Y�.B�"�2UC��\t�I�U�7 ��9�7Gu[9�p ��xb�C���g'koL$Ă��L'�4��A��C�4���c�y�52"n�r��PXX��"���^�r몙�sQ���k�W����ؑ�ȁ�{wj�@��^:&� ��4�f4�{C��{o`
U�z*6���m��xn���  Z��q�pb27A�D?���i~�nN�kis��(ġ�8Y�7������ܦ��YN`s!m,��{�×ͮ{�ZB[&���T~���e��T�GB&�wJ-Q��-x	eQ�	o:y�-��˚.�{�PJ%��L.C���ɮQ��Y�@ws�ɫ,�o/s��ݏ��O����t���'V'5��<G�r�[�R�X�tlkX`D��\|�p�T:9��Уд�����^�����T_~���}�M�#���H�$|���,y�6kNl�7���]��X=�}g��t�T�¾ɯ���f��x���@\F]נ���I&������1'߽x|-��+GXG&�hj���6:ӷ|l�kBs�$�ς�_l��-N����9�g�J=�V��|{^�T�!/66N�-��x%ǡ�q
ɍ͌h,�ߖ��J
�T��VP���w������З�"��:kT4 OQ�ߙ�a��[Q.ڮi(^����qv=��"��w����=j��P�M-�=�<E�9�S���Z�F	qmX����b�ԄL�׾%P$~�%����X�w̸g��#�+�/� \�����<�OπbJY�$�h���'���N{lP6E �B���ϰi}��I/C[��m"�X�$e�N���1}�_�.}���3r��_���j�G�p��[�p�L���&9;֛�+_	����/s_� &�����BC��LH���ȥ7��U��jl��;��Q|-\2����ǷEc��]���m��ks�;�h[�$���z���D$�,�^���z��H�S�=rݚ7)�`���
�O��Qڂ��>�ڷ@�$�/:f���qU�m�CSpA�i���ߢE�u����t�!�i�B������&)�������C�Ɍ���C�Wgv����~��W�m��n�lF�B����"y���@o��;Jy���s�}N)��]Ib���&mf�(o�5\F��"� ��/�5K�<���+��տ�9x�����D�����C� S�쓚 �s��(�*�`O��e��ɩl�������^|� �2p�"���\�C����հ���tP�РG܁F�7[�������Sf�����E:�V6,���z��Խ�Ca�6qN(T�+ё;w�GڛjE=�r6`U���]�QO�C��ӵ#�m���� H%]�@�S`�s!,��
���ou�Y�려-E�5Ǹ���0ۈ�C�Z�[��,t�e�E	p��[�k�e������׵��� �����HrF��<��_�^�)���:�5�	�΃��������l�ٲ51��M�2 {;�t��@���ԌʂRR�[�G���X𨈁��d\θ4��#���f�a���C��Űz�1�&�w���bU����Iyt�N�gP9��[�^}��,HL6Խ�3F�	dx��2���-�GC\}�����d�%�j\��>u2�Zc���V�"���w�@я���)���V��i��l�A[[==�h;��raz*Uwi�r.���!֌��n	@��"9��4<I��r�����6o�k*�3#�8��	ݮ�}��vs����2��DA͐f�@�4e��~c0��t\�_���N�/OYc�fi���T@�<%�t1H��}�����H��pPȰ�\���B+?�\��J�ͱOp\V�5ڟ1�zo&�o�V?�����DM���umL�dN�llv�d��u��E�q��,��k�n��D$��b�ҦpE^1��\,4X�N��D�ȔQ��� �C�����Z<j&f�����^J�h4"p����*g�V!�¤��w��3e�9�= (��>R�"fwq%y�� �W%�>K0��Cvr�%�)��$�wP�>������p�1�@)i��m�8-�^5h���gj�C�uF��B^$>��r'҅�K��;��:<�|u�Y�>q]�u��C?����Y�"j��_�?z��L�w'4��"`��K��.���a�G�Q ��ƽv�j˄A�}�|�r��"��7P��e	�أ�}��N����z�������)�`�1}����9K	�)Ч����?j�۠N	�F�$�K�f`1>�-���݉�?��c'�o't;箓h/}��-���Yc�eH�ϰ_MDѾ�� ����,9���ǚ�8VdOx�����@Na����O��oM��a���)2ȯ	3�i�>�.�O;�����L��b�D���K֫+�!h'㇬���M��ٺ�4Q�{��2�4��0�_"N�v�i���ȫ%�u�ͽ��ȧ߂g�E�����:[�g�t�M
����j{'��S�8oP��Ǘ��&�9���ߜ02�K���4��(�}�Xܹo`�J���r-m���7d�NZ)�/4��2Vu�8��9��F��t�X7�^8B����:���(P-���h�y��6�;)T�!E�*>2����WᄂB��p���NkSQ�gˇJ$È#���	!w��'D�� ���Z.�O#ҋ��̐�˞(�K�X�Sf�*��B�7�V3%������Z~�[�]:W{zj�#F.C>j��<��h7��
a�l#���4u��,7n0�~�;����t�;����ǿU�q�Q���[�b�3���<��k�(z�Z��v?N\�ԜI�>*��tB�k�4"U���"��p'h�Z�ι�)6�>3!N;���
�:%1�?�i܎����J�u�P���[�ո�m&79���	Z|Z��+��&A^��F{�/|*	�V���--x��wS�E]o|*9 ���Q��/:��$pq'o�i�V��F�+:���ch��H���hє����۱�=�׋��� ���U��f��}[��$}�Io~mqC���o����!�}G�G������ҧE`	\Λ�Ư�9�c�wG�C��duH�y�N+��gy_��6��8/��|�s�����esHԔ�&����.	>��T��G�q1�Oi�i��8x�竑�e��c<8W�l�����K~sw���R9
t���~n\SzO�k�hH�R�ʥI^��:SC�ҕ�����'�τ�.Nq��n%��ϮX��`H��Y�:Q�{:h �D��`�/?�K�<��,o�*i7D'y4��h;������1?�D�A�l�<��v�B6�ߒ�Q�<�{4�4ޔ� ;�i9W(����/��ˣ����AoZ�n;(����q�3_hRL��iRAEĺY��t�Ԯ�m�2$4�2i)k��U�!�]E�!R�;��Ht��w�;EG��[�uFN�dB:�?��0B˥���U��q���?��Bw#���5�QFs\�K��D�`�и[͝�My)e�炄�{����`���w��� L�>�'�$%v��q�����L��;5��u�]XT����_MGWu���%�8�#f�y�� 𶣹F�TvBq�:�l�m@I��ƚJ=�=�&�����{��Yz�p���(��̨�v��%>
���$K"�>�������%�6/h�*�6�塓7��Ƙ�ًjv�^���[5��?�i�y\~�Z%��l�� AD�������Fk1RR�w=r�F@ƃ����/Ȓ-�i�MA��?��t�b�ǂ"�X�-:P�qJ���M�U)�����{��>���0�o��X�m��HbZ&>�oq4��Y�=����R1�qǝXya��0��`����5ܦ	v�ܴM����ɞb\rC���\~�#b���a�G��Xw��d45���!+�z�jі���O�� �ț���ar�m"Y,KҚ����k	JK��;��I��|�.7�e��x��┇��wo=	_v�	%�u&�I�6�=Dcd�t	_?��?��z�v}���!R��0�a)U<�|�oc�?�HT��M���Z��J�۫��1���t5o��g҈8�����y6�lӠ�� p}�ȳ��3����N
��A�ů^�3}�`�c�H;�aP�$����]���)�K]\Ո)1�sc�֥��P��P�����?�a�ѣb�1/u[ �
�������7�.��Mz��ß�1@����$C#�_����4�ׄ6���V���Bl�q�hE�P猁P��c\�-!)*����~�]#�`��*��7A�=v��'[m�?��Z
�������)?�g�'o3�K3��c@m2��8t<U�L����
��}|��2��6�v "�x�P��X�"�!s0����3e�U��(�����X7�A�.��z�i̯9�inUJ��s8/u���j��p;�?����g}!X��o�"X�qk����d�O���s�v���X˸ֲ'^Mv�Y<�:BA��b�=Ņ�c�1H��I�6C,��8w�"�)�>)*��b�z�g�}�ю�;�)D��Jࣚ����=�˪D��ci#�	1>�]�s���y /�r����&I��R���g��!��EW䓲����p>H���� �|j6� �:'jI�4��έ��c�\F=�f��L���Rqp�s�k�@�4Q!��a��b��	��zQt1�h�?��,��BB���X�Z�����H�G9�iUv��R5�l���|J~ՋU��'4 R��B��Q�|>���NK�@�gJ�o�(�����BM�!�^�?����g������u�*ʿ����\p[�v����ji�����hW�;)sw���1
<�������	ZQVK�
s���Z�9��52H$G���%�H�G���&_}[v�R4��;�Ow�c��:A~��JkF��@�������tA���p$W�ʈс�#�հ�+8��9������Dl�ʟ���w�eD�0%2.>�k�a�v��g�kj�݃�;ft���	jb���J�I~q�+r�T72�d��{BG������<6v��9�L+iW�KK�)b&�� �莓]|�]�>my&".���<�\�	�TK������'@bc�*��������OU	����*�����l����;�A��1�Ϳ�G+cƙ������4K" M\;i!������%_t�ǰrU�g;��V��2�2�J�%߬_V{��m��3c�s��%|B�Ŧ�K4�M�='��K6k��K,��ò���Ir��4�$m�`��lp��0�5Tެ�:F[g&��s�fJ�����	��^��/O�'XB��eL�ڶ�O|�er�Y3�<TOc7W�V4�P���ަz����Ay��Dջ����$�ڹCb�|��l�9��b�b�������S"w�a\���Ξ��iY��?�0�"6�U�Y��$��$�n�&h@�н:���E+����#��&X㐊(2��z��:S�/hu슗Jy��u�o�et�+�Ӣ>��Ƣ����<�̆}U��`|4,���F�JtT�����#��Mn�a�_�������k��[۫��@p�h�v��6W�XBi�p���W�"�3!?��q!L��)�

�k��0����Cت���!o#Q:N�W��6�%���U�4�:M�3zI�8f��MJ��!�`�L�+4a��Ƴ��h0Q�dBן�^Y%gOC!S���aSW����/�x\j�/l��)ui�o�95�|�yׇt����Mjo�G������rRa��@̓���DG}Pɰ
�z�Ylv�c��<cl3�ZF��v��RKr��2ݹ�װ���1�W��O�(��_֞�M�d���x�zI�8{ћ�ћd�0� �+�dv
p��|�fͿ���	\�g_5���>}�1�=2��"X�����>�i��S2^��ŧ���`�H��߫���ъ�� �KSy9��ŋ�Cq B���Xy�_�a=�q�,��`*w\{���P[��5I|gȰ�O<yA��c!>�V��%�p�L�]�L��X��@��R^�ކ[ nI���]d?��;��1A�6�{>�֜�ۇwV��omsU|�4��2j��y5C��FJ���y/5v`� �q�}@�5�׿2N��/�rByڠ�j�S����$N�:��;���J	�޳#Hls��(��C"`��#��R�V�\z6�ؽ��*��Kw�vKt�7���ZSQ���Z��E��I��W��O�_��+$ ,=�I����0�[o͝㸩����"_�_(�9�Kn�I-z�b��cb9yP��L��E��s�����}�%b|�������z7�	�e���;U���Q�m���w�gr�qb���d�N+ف�`��Z������0��~����ޛ��6�3kkf���8;!�s~m�p�HG`��16*�-�5�ӏ�' W��n̑k� ��_|0��n^r�����ڜ]���� �^�[Ip��_�:S44K�\7�x�~�PD$2�i��oa�%x�|9iI*��q�r �)g&�O��\Fȵ4��è*N�Q$����(�PH?�د�Oݏm龟�h�>v�MDIb>�0�'k���à��γ��^hb�+|�F�іUv�m���!7'>,�ܦ>ȹi.�Z�b8H��b[ŧV�z��'��.\�.�� Yޖsmo�<�DB�
i�;�'�˺?�2$w��=����餇��wR��J��k.LZ��o.�6�?�C	,�.�࠭� �B"�/7��T���|�oY
����M�K6}��n���X;�{��?� 89����\�vI�l*ᮨ�rj׍"��U�랈�/��_��ZD<Y�p2�e��aqD�>u��0�MV��9�!�u����R<9�|,�w�� ��~�J����<��^�=y�Ô�,���ʒ8��L�8����GԒ���Th����Ga�
��lJ�;��N3�e��)�=Q�U�5�˦���{g��J,���J�I~���{�f�ͽK��D!H� RK��z�5�����&�3��K�T$r: �M��X8�jF�q�} �cQZ��A�{6N1����F'͌+$�<�4+�>��v��bⱟ�0kSv|*����e�p��Im�FK��^�r��8���A�j}I�"eH)��D� ��bQ�L���AgS|�$0�-ˆ"QX�p�Qq|���{|vB+��͝�	��,�L�#OI�b̲����)Fb��{��X�xpH7��d�w¼�;ѯc���.�@��h��}*d;ۯ�G�����Y��?�켼� �J��}��/1o��Mu��"ѷD
5�Q���$i�uǄ2�i����a����}����++�mjɄnW�6d3���m�ϊ�����g�.�Q�ҧ��K�=�E쀪�Οl~iq�7�ip̘����w5TUo�ٙ�)Q����#�A����K�F�G�8�ɢڔ�P�$���T�ͅ�v�"�w����D�&t���7�Rj�_X��>>Y+�0�G��H��rfdV�W[Έ�m�I`JY�f�2;>l�Y�3�*��j�d@k��ZH)���*8X[b�?ﵤ�
Xh������Ģ�ξrq�3��m`�S����b��Z��i�� xR��:X�U�Vq�˻�5Lծ��K	�b�N����e����`�Ԝ>��D���J�=��[��/c��%�l��H��;��&y��:�
o���-������t�[�8����� ��K��C��u�.*��"��8EPcJ>�������T�BFx������R2�O,�,�ͪ[�}�qD�={�T�\�u���=vj�m�1�X$jO�\[K��_�����c����P.3�X���C�/Y��h^@n���R�q)�K:, z�r��ٽT��ŭ�>	�$<��qfS`�$T��&k��uk����=��M7{;m���c�abGv���zKa�����׭�b���jV���_K���-����0�Z�բ���T�E�^~R�q� ��룣�9 �޹1�Pb-�' }�H�i�`�Ǻ�J�^a<U-����L��ͺ=�>��y�.�S*���x�����ЇDdi�d];ITG�hv���;�+g"C2��cNylJJ�;Ks����FO�`�L����Q��+����(���be$���Q�6�L7�jD�~��gt�k܋����AQs��^0��JU{,��uE���xA=\~���p�� �����>db�М�+�a��l/t���!���QhOx!�J�bs԰<�d闾�:g�C6��'hC�KV �����U�){�*$�'E�A:w��cx�Δ�W�{׫L�[�/g��&����|o
F:��[�K��N_Zh��.if��Y�N��B�h`7��ڜ���W�ي�����,���N�^,SF���=z�#���I#�_f17Ņe{��~z2_(���$fU��%`& l��x��>��rn�7� �ێq��h&��PH;Z߀��.�W'��qb%*h�G��OA�U��&�2ğ�*�-���"I���f1�G�?s-���垔�Ϝ�(�4%D����-]�����\~�~�1�O�^$����I&�\���u�K�c��7L1.��(z$�N'"9k�`�&����歅jE�P�\p"8�0�!��r�e{� .��
(#߯aU?B��=���.��fw��]bRWt}c�	���о up��{�?�G| ����fxJ�3JCi7bJ��/�Giv�:�������r��&�f���7b�Y�{����<(�a�0	9'8�RH؃Az��$9&6p�(RM-(�����X� ~�;��Сt�"�S90�~@ďjX�B���;���b-�@?Xt�6��O��b��i��q�@��_m��L�2Ks�H9�X��}2�.Zhm;)N��]���@R!�����#w�^K{�'b����Ŀ��Z��%P+�oq7]ιQ��6����E!g<�%�� �Is����.#�c1�B��%}~u|��ыL�\�I*f���{~nlL�.�A��I��Rh�V����7�p6ve=�����"� �C�ϫr^,�G��MՎ�r�u�ܾ�>�c�̀mAd�._�Ш��-�g�^��PC*F��{h�x�x6�A��r$g�/��F�a�<�Nb��/��Vg�۹�lgǗH$�"��"�$Ӧ��SD�3�ũ�Ƶ��{,��l�����COk��4�+���-O_/�xI���:�_M��4:�$�R�7�GjQ�����O����U�{e�iX�	�����=���pe�|b�5��\1����t�9�|=\�8��^S"^��k憫w�o�4²Xm(��o1�=���ץϨ=�|����g��k��NȪb��|�A��C�{lB���5Cq
f\���7e܎o��e_t5���#���P��q�QF7��ERP�<&�l~w�˵.��!�j��^'�MUv���9٠���dC��%��?^�t6@o&��D�>
D�ZH���@[�2�G��"5_��<����r֯�»�s�o��'�ݙ&6󶹢�x
�ͦ7�r�f���:"皰��z��·��F*>T�;͉aʱcOy�8nϩ�M#� �����<�g)#l.��ƶ��U�G�=� 9�9�E��I^�A�S&l��H���[��`�)�ٸ\�8���q�s�Z�	�L�:O�b��C�iK�\����P�qO	}t��Wp��RTF3�-�:��j�Ͽ�jS&K�g�q	f=L�&L{<w<���$SЯNv��j�d�m��d�������&�T,�j}�mM2Rţ�?��S�x.���X_���ԇ�g���ۏ������}B�'$�?�km����d) E���qұ�t�)��E{	��B9�ߐ2�x�bȇ��=�4>�#!}�+j��]�����zo���v	�q�d*l���˧�wlo���IELu��#s}�[��XO�E�V¶�j8�j+��9U�ѿ	Kc�I+�]{DH1���	��#ʳ��)��˗�_-�W�N\�pCSM�_+Z.�у������dz�í���2�c`:uc�M���	�D�G�h�oS�y�ף���Y���lP]vǃA��}��+�$��N����ޭ�w���X��nfU��QY��!�l�ݽ�Y�.����t�����2�m-+�ɋ"�DhKU���#}�´�xV��ц���>�::���R��5�;�U�����)��d�<�(�c�C� �h��=6~�M�VRxzڬ���р�҅YGf����\��p�B��[7_�d�T+�$v^r%mI`���X�J�$����:ˣ��i/���:�V���w�U� �A�����pf�O���@\n���*D������Shhڗ�F���tl r�����T;��J��4#�*�ǯz���:�3c�-�$�]x')��ğ�|�f��vbs��ҙ����^�e�����f(�;���hI��{� ��� \%z�RW�X�'s�4��&&���d2T�fhv���b���D� ���z�:��)#��^s��v�c�$U�Х��#��59�,Y\�O��P �R X5��÷�{8��'w[�/�>�/�6!���/Ւ𣣟xp4 ��sl2p/����ߧ�{&���;�>@���h���#����>�t<�;j-��}����I�U�C�{�s='.1����� - ��U틲q�Ҥ�'�I��K��t�Df3 \�֓���~�H�z7k���j�V��^�У����G���cDxn���  ����7���[�6+��Aa�Ž�;�D��L��Y���=�ӅL�)�ܾc�M�й�����.�ԧ*�S1��&9VW<N��R2��SIM%�%�a\��e��xs��`�K������ۓ�׫y��}�&�Kd���+�/L\e�t��j�#��͹׼�)C�F������=�ꥴC��� %.�KJ�g!]6���tQy^%������:�h	\l�eWL�������
���~����a�1�`&��b�I�z�b�e�)a��8颷�������A�L|IƼc�1�H�Ɯ��_�.����W��� u��F���ĦA]>���碑���	�r�YI�z�t�@H/z�	2.�SZ�L�\�u�I�:��<�=v31"�<qR��$��Sc��
���8�����f���V`l�'y��A4��XoF�ߚ�X�v0��mt����ۈ��̥jU��D����d�"��ҍ�����ި�#�6�>��}�/h�af(�IӪ�e1b�P'C�n�6�� c!�c���@u!��s���+gHOO9`>b�s+(�2NW��r�����0&ޖ��6���#��������fEeK"�҇䚴�_��WV�Z)�pFɞ������	���HW��������R���E�mP�"j?��.��u�f�V�0聼�o�<|R�?MFj���ڎ�x'`̢��7*Ru𞩭~>Vz�I���滤j�?�Qp՘����5dgz61H�(y�W �RR���ch�S&`�������6��,�Mo7��ٱ�w���w&��3z��Hh玾��]�&���9��+ާ��˸l���E�Y�1%^
K��8l�(���W�G����V+�ܚ�QvC�ޕC��_���k6ܔ9,FQ�~���v"3`���>]P)�qg�{�9�*�Po��4���
�ȝ�Dz����o���?!)5T���/���#��>�	�$QWG�.�ʑd�֣���U����kO-5U��;��>L��6������+b�χ���� F+�r��G�t�k;����+�
���R*����!�ǅ�l�$�����L�����MQ�:f��VX���������L��7���<��T#V����-,�˺��	�=����~�)����x�X���������C�y)�G�Y�=q:�UY$�8�7�U���G�<��Rk�o2S�@Ӯ{�	E�舥Vc��K(�#�v4����G9��6�_�`Obܐ��]�]Ea�bL/eD�o#�r�LzO�gf�ڊ�Y+�a��C�U�+���U�2E��R�jzz4I�������������Q�*��Lo��	�^�Z�Po��$g̵e���y�h�Wb��&����7J ������j1���n�ό�- �c�q�֛�g�l1cUV�^�FR2���\��3c�vZJ���"��2x�ԺMyZ��a�8'l�V��̩2!jW�2�W�o�E�Fr�{Fзd�}N�#�UΓԽ���I�����6�ݞ���D.�$g�$�l�O]����3սEk$�ζ�i�� v��M�;��34?�S����^��Y��b!oF;l��Y0��0�B�a����6b��Z�yQw/�7���Wy�~�u0�u{����y�6�F������s�ww��Ivgb��Z�Ț��7V���J�ܔfC�|(3��ݢ��2�`��J��LNi��8e-��)4��;�U�׿�JaH�#�q|��"�k��A�m
l�Wɶ1�����Z�<�4����#��Z�0J�E��u�"�)WN��0݁3�R^�r�L��D�v�,�O�]��_,|�T	�1o�1w�� _/��L����>v�����<\��^�e)�/.���߯$y�*�&�NО˫��q�?m�q��o���)�Ğ7[��˸��d��gb����8�ܥ՚��vY8I}���p_ۃQih�c9#Bn`CĞ�����1'�8O��;�p�� �2y��mi�R��/�H����H�:����i[<�jqX��lƊ�~m #�i��A�������Ҷ��F b��ʇ�s:��^��t�l��O7i�ZFh4��l��O��/�@�$F	��XI�_���[�8m>���l�뻘!�j|�� nL�Aȥ�l=�C'�B��+B��ь��a�h>A(Qc��}@U��Ǔir�l�/����y��Z���%l�ႍ���`�8Rp�j���  �E����D
a�1h�ŋ���tK��|q&���f��P��E9���O��ӳ:	��ڌ�n��h-0D�"�
���T�Eƛ���M�4�dJ|o��7�¶�����e�4h@窍�.&tl3L=ɦ��L�綠xo�Mf�F��9�5��#�m��@����c�a�,RZA�~|� u|��Ѭ�D�m��28E�آ? ���J��H��Jj�|�=���l�	G%����8����	����E��6�.�[q�՛�PP䘿s���l����z�пr�C}������\��$DZ7�#���~k�K�������_r�	o�ن�]�y���S'�>>�0����5I9�yֳŤ4iq\!�ShĮO����� �ؙzЂy�/�#�o�1�:RO�K�w�������eQn��js-��<2�o�%�K�ހ��T[�#��V�D��� �f�ce[�M�e� ቺ��_R0>0�9Q��U��G�����$�pmY����	��_T�}Q�}�}�he�r�􎾬�b.�n��,ŝ�D�됍0�(�,����t���3�K9��ڣ�����}�܊U[P���^�|������;����0k!m�5��h�w*L�:�OP�2rk,(eL�	�a�����P'a���/��������7�F�ךItv��%���G����i��Zj�#Xb�)�7���	j*��$��bY��gv$p�����0D[����`��"���!R�M�\�#�����l�O.G��~����ԔJ�GаR�T�54�1>?3�����ځL=��G
a����5c��|����8|G��Jڪԉ�O�|�B8`6��$ }	�L�<~gU�\+u.U>\�x���:��/<����J%xR�	2ep�"f�U�}Ɖ�):D�u.ߤ0%�Y����TI%��i$�>58�39�ŀ<^o�@H�U�0�����W\z�9�`��έb=�qI��v���OrW���է��5Ly4k%8*��{8 _��8-%m)�*��V�R������t`K{_q�o~��V����'!*��t��4߿���,��"gR�\����IA�%��l2�����Φ�D��i�?�kD(m�z�Uj�e�l��ʞ��,�������+����gC�R���`V�K��֠�ڥO�Zc��@��uW��{h��l��+�t�J�H���4:l�ر���f��كe��=q���dU�w�б�o�����}�	ġ��ѽ
Ϙ�r���:l��Ol�Q�gq�� I�F1s�+D����`��(�nZ�
��U���)������=�h:t��ƒ�2\�-*>9#�v%sմ��E�V�i��jjbTwܸv|��[ڽ�.�4��֙���#󠵮���Ít�P*=�䏼���������Q�$���;�o���B�ӹ���^k�i���8MF��{�%��'�L��WUP���zr�)ms{��&���${Ǉ& ��4����E<_L�*~�q�!�]�%�2���b3sc�yRE��L"1$M BhT�e�b1��@���������]�xdpG	�e1>m�d�"bW�r�`�y�D=y}/�}�b��"���z!�}L�s�]��A,����4���$HI�|Z}�|.�%��Ѓo�`E�J���X����|��f�
@E�^o���p�h*�a ��ᬙ^_�X�ߋ������ƕ�Nn�(s
����S��6r�Mq��*Ӌ�r�_��+�z���M�Uc�0���9V��Nbp�I�w��B�rj��� +����ߵ=�౪vh�|���e�	���Ɛ^��A1C�eT�b����a����@�Y]���=�\Y���P��..�4f������,�����}��B|� k!�{�6	��h9�N?JO馅�ٝ�u�a�� �d^-:5?��2�7ᩚĶ��������qPrv�g���9��̬F�c6�u�^>{�'��_�G���9Pk��X�� ��e�:j�m x��XUĤ�gK��h� ��g{A����"U��a]��!��L.Y�U����]�L�v�5g�%��.��Ŕ�E����"TCH�oFV^���ٗ�e���-[����O�4�A���y1/�T��s��$�y��@�"z<��{=���G��W?�@a���J3�
���v4��G�]�,xm��qz:h~���3�Z2~�X��Z�R�KԮf��9'�CK�y�󘏮������o��1#��Hb�O�Q�.	{���Z�Θ
z�:R/aV2g
1�!-�b9�X~��/o��7�E�ߪ鹨�&�l ����Z�(�yX��_�U�!!��"�p�S�����d����{4']�j�Z�h�';�����s��"�2���G�U(tK�;�I�D�ȝΈXUӖ�h�=�VVu�f}49[Ío���!���p���$��͇����r�FnU����l�;Y$ ��>��av<!�`�[n~�\�yu���D���_�s$�GZ6�깥R���� ��
�i9�*닧|J������{1h-N�_���_q�'�6�s/2���,5j��+��zڊMw 
M���R�ts��<��|��MP���ͪv�����Z����7*X�6Z�a�V4	��|���19��2nI	A!�����]w�h��l9Y|��W�9�oR���h����)�?�õ�y[$J�U.�n�Y�'L�̎�R�v*���F|�O��&��4j�{�,~��I��	靅�?�� ��~���՜���'�1��o+��P�Q�W�;Y�e��#���D���ǖ���1`��\;i�*gfB�`�S���0d�Y�Ƨ�M)t��y�H}���\nF�6�@��Hu\܊F-���;mpvN%E�L�n�=d���ԃ<��<ԕp!�����K|�l��N+W�ye�4^�	\�?4���ɖ?�v7�%���fX��c{R���j���-���>��u���l��=Ŕ`�`���=5s��P��\:c�R�ހ�$��x���Fm@3#�qa�U��)�B?X'�V+oT~�F�Sx>n;:C��hu1��&��)0D [��A2��NN���p��D�� x�!���w�0dy)�r`�9�-*7<�]'�Oyb[u]��G',�V��mpsѧr�mOB�tO�
�x����U�җ;0�1�V�a��*���3M �V��oj*׼�׎�f��^�K�8����mj��c�S-ԏЃ(ݴ#1�U}^G)��ݨ�������28
���ܰ~�s������iR"�$��&Cz�3ŇR�9�+*�X���}	�A��p���w�n2ɽ]���(�9��v~V�֥E���'|�S��gU��Eb��;�6M�Yb��y�]v�R�~`�5�G͉��L
��h<2Υݼ4�{��GF�K|s�cWּ�]�Pm����xN��=y�Hb�e����E���,n"b�KT(]�`ȥ[�
pm����oF*`�>�2�g'c1��*[�}|:��]d`{��,�վ�	��A���L��:C8%x�9�����SsH44��cj�y>�m]�ԛB��������6���I9�r��<���N�{j���<����%Q���%J��iC�8�U'�V��J��a�b���L]����������:��x̠�8?��ϨM��dDJC�j�yaX�A/0X�@m.��Qy�����bW���AR}gr��]f��͊m�W��ݪ������<ϵ�(��!����Yr>�}�����5 ��1�W��zO���(\��C�����%O٫٪�z�Ne���,J�,qcպ�YdV) ����t��J<��H�L)�����}�#������Ո���%:�x-������f��H�1gX2Ϸz�?��~NA�L��U$;������-�!�ד���p��OjX���O{�b�t8l�DT}���~������sv�2�������I��f<$�B�l��0�V�]��NQ����>Q}�C��"�I���f��M��{4q3�Y���[�����T��i��=�jJ�.fῂ���t!E��{�V��:7�fj�.��pw9�(
Pg�W5��u��M��X�m��Ke�@8-����o�Eb�[N ¹O�*��03��|L*٥�&C�5������]��\�Nڜ��k~$�͏���:�����sjH$h��P�-�)�$2�^�l!�	�w�z���7�
yq��EoԆ��ؚ�nwTOe(I��"t�dx}�'V��}xٛ�7���V����/�O��G�2���΁���̴�k�.���W����r���.e���C%����u�5����:(u4keB�����^�-1UD�&P�O�
qCL�u�B�#O�`��3f[���������I��pce��[�HͲL�*�D��ڹ���cʔX��">� �(vVs��Uq���XL�A���h��`�ni)L���H��Q�g�Pm�Tz�o�j	v��勾��G	��-^N��9}��=v1��*�a����d
���H��ٖ��g���[����o8��~���밧��lQ9�~"�� �T2��y���(�{|�8�&
Ǥ ��{=m�l����D#E�\t{�Y��LCqzUg���:͐��H�5�a�n�7��o\���>�E��e���0�H5���ya��+�2���9��,����uznh$7I}�f�٧��&<�dU�f���F��G��_�{cNr��6���a�I�[Cm[,:�D"�V�p�����7x)�g_�砉o��k2{0��,���y�jb��7V�i��_�w�lb��ȼD}������p��	J� 	���w����`��볡7>�.ވn��O�I�*�FB�S?*7��H�)��V<p콿�շ!������ ��<N�`v&P@��`��k��V<�{�-�k_��&�Ψ���ڮ
@�ڢ�O�M���]�|Y�W+m��kDT��r���e v�␪�kh7Լ����ס�O�(၏tÙ�b��\���Zl�_���fj�h����0F�:"J�_��}r��7���������yp�K���� G�P��2;�y�s�r8�$EA��1}��Dp�e_/Ϭ8�C���	����R�u��^z����i�[�KՆx������	�sQ��-;�6��S���h��fCD�Ʊmtz�Č�f{���KKm��(�v1!��0��<��'O� xJ+���v�a�,%�̒��T9�L��|βƛ�t�x���%���Z��l�K�颇�tZ�2y	9���-	�G��-��P���cg/�Mj���'n�����l*Aq
Lp2�(H!���g�hBX���q���%:�0P�ȮE3*g��☃"X�͡��Aos�v��U��8�o�����r�����Ҟ�!����m��&���A����75b\0�~��"���_v ��^��,��ZKi0�upy̹�� ਌�D�������>n�;O��Ѽ\*��p��AY5��o�C��p��v�{ǒr�ѥ��H��`ʊ�5u�&#!�q��˼�u?�	j�Z'7n�퇯�Rxn����0��!�<���2V�o[��F��~�U�Sw���Eڊ:��T�a�������Z��:�=!�'�T�Qe���B����<"������*���W�p��)?ֶ㥦�7��}�Y&vF~�"(?�VmwX��d|���)�W��C�K�qER��	V������	x� �`�>(�������
uG.��s�_�1��>�R��"��Ǩ������M�^۔>ߛz&,މ{+��R��c�-�Hw�z
�H����a"���+ՊB���V������Rh��-��1�AO~�U�wC� �L��lVJE0l�E��	N"\�^�����a|^nY��Cv^�6�j_ ���mQ4�ͤ�̷(��������%�n,�zVp|B�3)�H*�
��E:���N�>2M��4*݀�EJ��/M/u~=ʓ��d�*��g~�׏�ES�����C��Q�T�z޴�,-��2���0�a��`]�qq$�h9���U0rp�o^O�6�x�M����'��l_�X��t7�;���來B<9��j�#�K���ǉ��)�T��l�`Tx�{����+W�ͳ�fHgdUL�`;��.�d�g��bh�A�e�7ۅ��6b�.�� ���f���[���\��`G�Ɯ��?B�U�w����k�A�;��3M\j��/m�ڮ�:z}�N��a���9����7~A�C,����}�[W�}+����
��9k���Sk�y1�_;����aRIcA(�X1X����;�=�8V�ҝ�"F)��� qlQ
��J���G�]7x�~�a�-s"b-�����vPH��/�No�}��@o��>�
iE[��d�p�d����l�\<��5�K7;����fDj4 1��G�W
��C4]��E\g�z�:P�T���Mc2��AT�U�s�U�Qљ�;=z�}�8b(�/2�Ѻ����8T�qgD��C��Kgv!�X�bY�~�z�-W����3[L��t�.�Onł�Ӽbb� ���B-p2�����~r��G�z���e�X�=߃_�RfA��$.�8��:�}��n� 񓊗��)��h}8
,����%������M��Yµ7��S|͗M�������4z���-�`�WZ�q��*4�Y���M�Nu�ע�3CU:�xJ���մ�իF<�����wC�����G�\�l8���Ъ�_��j9Э�[������ƀ\��6+�okv��{�`[ݖa�"%g�'�2�R����A�� ���(Hr�|��v)W�6��0RX�".ēoF����1qs�dW���LN�imV݊�����1�Y�p0�C�㼟Y{��}�����������UQ���<'�SpA��O�2i�̀:��l��%w��
B��^A���t4ϕ 됥3D���u�|�W��/娞���g�+����E�"���x?����Έx`�f=�WZ����f|Y1,�1��t���Q_VikmJ��S�c����Ƈn��`�����n�9���)�Μ0�8�-��P�O�S��dX���53hr�i�����T��zg���D�}\�e�V�b�5�2E�Wrx������"E���������E#�4���#S�th��!���F���~TqJ1�HQ��}F^�|��0)�HCu�Bwo}��9�M+��z[��H��(aR�	��g?��ԛ{Aju)�_F+�@��ɦ��Z�9C:��6�9����,Z�(��ω���I%d�+�Q�675�/����3q���R�Om.���C��o.��9=଺9�~��b,DT����>X�i�5�K���K�DLS��'i�d,N���f'8wz�qHL���KU��� 45H�����]�z���8(��B�S=���廜�̥�g9�h��pT�)�y �wb.�Ȑ��XDe�7X4�1��ֺ̈���6�� �������SE8��P�����t���zK=7��x��)�����m���7{����Z�E��ǯ�\����:� �� �SǺKŒ����6P�2��笆��������N���wm�WP^�`�`d(�x-�uA����EH)�n���5�!��͐�4��W�H�x�v�:�������+I�	�r�e���Q�����nF�-����gg3����p3��s�m�lg���tӓ	���۫��2��@ϕ6ڲ �lS�����_m޴�7Re�ͨjx)R��U-�))� lAH? �R�(�I�3(����j�G�k8u�U۵;�5�q(�ᱚVb���3�T�q<9����b֖b�s��r��bDVyY�0�:@;���/,�rC-�u�߾�X)�F�h�q���Z����R���s��2� �ڝ�;���p�V�B��iR֟a�CY����R�ѯ7��8�9xoD�0�V�l���_�����ciH�7)ڭ�kX��" �}AU����ύW�q����~=�\:���Ƶ܂~�� R� �� �������@2�w=�m���3i>�p�����v�ދ߬~#��dյp��?9ˇ�>���0�Ӄl������3����M��I����:���P]������S�;A|��%A��,N9�OT���$Y�E���gs�vM�2	l�~ʜ����"\�{�`���xaSy������3-H���#�8n�=E� %��cWΩ��p^[���ǡl'^}k��I�xF��FH��W�� kw�CȁѥR,����êr�=c��YM��g��gװ�4B��M!�4w4͹���.��Q���6 �\N8�a���=��pO�D��'b�F%�������n��D��)n����pK�D�hf��Z��z�U<C\o>�fw���pXz|&�����;�p	벬�W��|��o��Hz��'�����i
D�3϶�bu&�����l�+���S)�ۜն�����<o�Bno+�PJ	-�Xh�ǟ!���F�<�����斎v�2����RK��z�Z �TZ�t����>�
�X��[�Uҥ�[E(�?���ɝ�i��\�������1b��#��,R!Uմ��d�<`��Ԉ�p&Q�g�|�=�� ����h��@қ��P������ �!�j�N�<�*����/�3�֜�R���|o�%�8d��OdV�=y��զj@�cu�^<�0n�ʅ�:�t���!O���.X7�T��V� Wj9R���I��Jx��u� ��>�>�d�f�)�:�r�<�;T&�ijzi�e�Ku$�l�1���e��R*������mo}	�n�������˙�����j����m)�nK�FO���'�$�mSn��-λ@>��(�nq������L�7į#�X%b�3��Jf�bR5���H�(�����+� S���ڛ�t=���/˥�v<�b'��GǱuM����4vȼ�e�3a����,�� ��h�Q3�Ǐ��M�p(�
������2�i��v[�BK�[U��ů%9/	,����hX��i���n],��H�L˄�+Y���I��QXJr�$Ie&57��i���V�����*���w�ܼ9���a����۞�5H�Ax������3�ю�=�1����A]�����5F�"��uE�x}����a^�*τ��{�2��
���n�d
5�o��������k��Ʊ��+L(�n�dO�wn���`9�ƌ������ę��z���~s*N�T�~;�VS&/8|�>�}�'z����-��2P�'��1)�#��ny��T4{S�L��7i�I �1 !����n7� L�{l\�?��В1�A��K���v�	�(�0��jȀ��Gg����;O�����_�W4\�K��X�ַ=H���U�DX��HBcO�[�0�G��vw�	�I��3J��AMV9�!bv�f��%*����c��xt��,7��y�x����Z���Ee�#����%�z�`b�^�QMMk�m���"�[X��-z��F#?|^��M8-�fB���/�+ ��w�H-�L 1�~s2��t�j�u��.��^G.�6���P������8y����qp�1�c��Q�G훈�$|F1��"8���4:{��D������d��n�A�m����$�׶%�$����&l(N[Ϯ���JY��a��0���'�0B����Y�����?��f 9ё�Y�BI/6_��p�\��P.[*����LT������*Qz��!yp"AJ��C���C(o��Px��7
�0
��|��#p�+�>P���p�2���jwH@�"F����{�`>,�����q��~�C�$��)��Ĥ�O��������p~��.ܖ\4�.�|��Xbq��"�߿Aѓ�%���)�����O�ɕ�'0$�l1w�Q��Խ�U��Z���RѳX6�� �>L/M�Z��/���D2��E�ʰ�K���2��pN�X���������=���S�|�-���^dc���)�?���G]i�IA����,�Qw���W!�����t��;#�T���\�5[&�etI�-v�7���1'�Pv��g��D�`e?���?�<�'��H�2�A�1��$����8O��wp?(����>0���<v�s�F��|���l.W3�6���𰒨)�:H4�u},����.�љ�х"���� :�(!0�Ҷ� �c�10;�H�3,�q����tLB,k�n�,Xf��*�@�zBs���������� 8�fL+��#�ⷢ�򶗚OtvO��ŸA�>���:�="k�_!������w�#�Mhy�ߕ�Bh�������F�d�k��R�6X3N�׋R#�6
��鑚ў) 1��=D^.N%-�-��q�I��
^,��P�S�!�)�tU��:�ꖵ��9K��r��V�C�=H2�Ck}�����V�0��ZS���u�����/,��a?����HB�:�[&I%/���LX�79�Tݎ�,�]%�]�25�@ װ�a�����n�B��g\��E2Co�GM3+-���]R��
c�qRk;ea�,�vK<R��*J�� �I:�Zl���FX�K��b8߀�b�(�a$f眰0��;�oP��h��·��`��l���܋�t5��BWp�����k�O�g1a�_$!��M�]��ǚfVd5�D���H�vD�])ɀl#��'��8�����(_)�#���"t��^t�a�V[׫�pڇ���2�#j����ߩ MB�x�T�sI��_0�^p�n,�jB ��M�@2����z�%�˩��-.��~�Tw�'�/�q�X}�iJ/z:Uǟ����['�Ry���� f����3�f��6�!Hr{��hd�������6����D��b1�tGi����a�V1��v:pq��o���/�5.;-
���^���Qv�^=X��jOȿ�7TV!fO|Do���5~$d���"/��9�?Y�+��n��DH�y�*��H���l����m�mA~��<J܀}����Vf7�*��g�6�<L,�BZШ��qI/Mun~���=Yw�əzrsM�ܟ?��DLy�������@�?H�m��*l��O#_��c*t�ә��l��ΐ����w�fc��߆�į�a>h7��/�9!E	
�M*��!�nghzTړ������4�R$Th��FEBk�w_���"+O�>]�MJ:�+��m��{D.�99�]��I��>WцK*����B�8s	[������6�۸e���x
���ݑHU�l�N��6�դYI�r�׏oI�'� ����C��S�R�%Τ�e�xo0z^IR����v��k���)�� I*z���	��M��o�@W�H]�;�X��i��e��o�'�z�B&	�O�w��Q����%ƤL����Z��󬾯��`V��=v��S5��D��^�5��Ϫ=�γ���D�f���%O�u�e\���/e��D݇tY���T�2z1;�xr����a�̪�+���e{�'l9m0b's.0����#�羪b*ݰ�D� ����uuƎ���_���0�T]�/��T-}m���I#+���Nk��^�n��F�RR=9����h��θ� p�1ZGV����]�D2��UL��fv�"b�{���
n���0[\$J��׶�m`������4Pg�O~��Y��y?E��1��&L)��.�o��<^L
�e8����K7��3��mΏC���sw{d�u��.�u��[|��r�����f-=����ɮEn�<l�1Y-��C�`���A��]�����&Te�L,Zb�[�܃�ڞ�V�>}�p�p�z���ׄ<�۪�Y:R��|�Y-r�_���@��姸&��vF�����m<����?�،��1_�I��f�Bg��T�`ɸ\&�!
 �_P3Pʖ��_>+�N (�T�2=�zB4��Ň�������z� ����b������1������ ,O�Ҳ<�(;�`�:�Gך�x�VW�:eS�r�o/�Q��T�����g�[>��EQ7��V1~�s��+h�%S n�V?XܔYz����>���	�'h�1-��>��@M��!(��ɋ�D��-�S�~O{��b��E�/$�2� ���2>�\Ea)VT���i9g��٘cTuJ�G1e�O@��8�2�H�	KZ�Au	�n�e�b�T��ͻҗ��yn�:[�?+��k�!�q��%p/.Vd �����UOJ����K@�+Q�@ �[�.{�Xo�U`� �i:m^V_/�w\�w���X�g'��6t����r�5\�Gٴ�Ue��e�M�n�6��km��IE�9
�
{c�l��#Q���9aT��f�@ww!�qh���AW˖�(�5�K�eD����B�����b>ְ�<������8'�$0o]��@O%��Ķ^�<M����Q�.E��죏w�(.��H� =�Y+�}�̉���M^�e��
oqL3���N�n��3�O���U��YÉ�R��I��q��_���*":�X_��a��ɂx��U��#D'&A��uu*ᛢ��`t��f@���b�Y��p�K�fF|.K�PBGqYInΩ�'J���h�w��n۱W�:��8������+��Q�C"�m��B�ܾ`�R��#~+2����l��a�!��3R� N.Z���K�N�Q׊ $vy��4���,$�0���saeGQ;U w1��\��B�&�H�Du}2I���!'��v�߈6�L+߭��+�2��~���=�D�T���M?��2�_���@����ƙ��otp���S)��`�v��\�O?��貽�`{4X<�⟿�ʸ?ͤ�'�N�-�A�%a�l�����*��s,nI�kf�m���(�~��'��[��k;��jU^6ڥ���d{�f4CW��*���Y<��x0W��L��X��~�Ɔ|�\�Q�%#\ Z��Pe�ء5�&[˗��7e������{Ӫ����k�bG��� E=�j�h�T�n.�8�`�97V�&��J4L��>'����.��sb��~=Ί�e�J�5���	X���v��w�v~Lr aS=L��f_�Y�!�X��=깁�^����~�md���*@�Y�fc���?Շę�a!�5B7vC���|�����%,�\Pɑ#3=�m����E�zA�Q�ʥK3��!?��[Ip�7K�BY�'��J��&���d�d���J��\L��'q ԥ�h ���(̼�E�
����Zw����1)�����d
6%�z6���40ə^��y?���<����uGI�*7eA1-HE�13.G���EhVa�q���Tk�^��U3���0Q��$~ ;���������6_Ւ�Ί=�����ٟ���(C��{�4m5�!U����ev��}��Pߴ�͚����Tt����(�Ұh��m7�[���3V7�S���R@G��F� =}M�t����}�iR-"�c<;2���8��'�x�i�/��u%	o�|ێ�W��c�2CGNQ������%��8'&+���R���[�tDwsK�O�s�b�I�ƶA��6|�m�[+9����7(|WO���(��!�u W����*	ڴ"T�BU{~��M����+��4�9���bZ��u��r�NQ%'Jr~�f��d0��f^		�g�{f��۫�����g�P����K�'\tf Е�>�L�a����<�G>}�!�i���DX�SPW��^�W��b�}������NNB���M����Z��w�my�7���{��a��k�&��͵(g[	y�����mT:986dG�.<S˿`i$�b� `F�lV�������)�K���uf�~|�޴���!?k�T_�T
V>�� -atc�iP`LV��J��v�����C������g0Z�%]F=ʚs-�����2G����)Yo��~�lX��>6���2��%�T�3(��.���~�<�K4E�$�Η0�B���u��s?��F�;��{�X�/���f3�I2�h�S�EnuNrؿ�jj,�o+PFրHw4]�T�_��V������:��;$4F����bP�D�5�	ZPn>��{���"� M��"��M9�'\���[$Q{��\=s��HV�F&Z��yY��+��̪-��%��z��\��p���IA|'!J���Ԝ�$��I��|�̘+�jUE�sι�*����kJ=Dh~?����<�m��@���オT�'�U�� )#?u�AΫlb8~����>��[�A�$=�8(�=m��J�T<b��3�ӌl��;-ݧ
��җE� H!��f��X ��hD֧Ř�	cl�י�r1��K{J�˯�8�@��} �g�"K�A�m����d����K#��'9�����@@&�t��RF>36�޶r[�L,��>�={��f���T�u���>��"���r.�$O�yhX�+�!}����D��u\�6g��j�����bS���,�����DV��D��LK����c��s|�����4R���1!?���^�Rj�!xc�N7�����gw=p(nځՕqe��-sW��䁺��-d����|K�O���P�4�,u��=x7�_�sN�$>i�j���H4�f���#�����BQT�V�ջ<���$H����PB96!vX)�8&*cQ6��SnM��B���/,^���3�R�s�z	�hB���;MFׄ�+�[������2���p�1���q����NN��CJ/,J���a8M�T��n0�`�X��X�KoH��-�� g��_�� !�
��B�rsCl�
){Ua׾,�Z�zSu� ĕM�{���I�F����#�H���L������L�WV���-	�C찅x�m��{�i�?U�漰)Ó? ��v��ɺ`�X�o�L�� �,0�ۨi3�:{ƍ)-:�Ԅ6e25��#^f�]2'�ݷ"����eu�A�M+�'ޱ�u�L׋��Ѥ�b(#�d0�4��ہZ�;��@.���W+Of����I��Mݵ��9#�[ȋ.DF�qh���`��w�O	/��ؕ7Z�z���6M��3���C�T�	Py�prD?t�U�T����xB�ɞj/j��jF62�Xy��"�btC0�Sĉ�c�Y*x�V�׺jf�J�m���e��a�`������s�+Y1�5C�k�7�DK/�/�{`����w<����-̀�>E�~�'.#[����CA�&�4�Aɣ���x�Fv�K?=�=���M�ig>WN%;���_Yi�����+UO\Hz����F��y�4��7����fȃ=H�:�N��S�� k���'r�9��M�r�x7m�Kz�ڹ(�� ���B
p1��re\�:�%�P�"~�U�Ȧo8��4;�lZ�6�aA7����e2��9q�S<�&�o*��y��6�$��
Ʃ��UuJ����/�3��v�?H�˼�����T���p�d7�+���v�BdgQ���+�4��n���:mVmh��+ܺ��Y��U�Öi͓i2��}E(`(2��Å���������jb�%��:���|���l��{�+mUd�v\'��Qp:�}e�
�0�g��I4����?4>���|�$��I��T�<0�Q3�h����5��S����D�[���:�w��?[���]ۦ �V�u"U��\�cgd���]H��O>�.���.�NF��c��gk�|0�m�c�pg��-��)����,�(�H\۱�r 6EP��ˈO����(p����ƞĺL���5Ҝ~I����̉�%qn{4w~�ؽ����z=`�P��+�؃x����*=}��~VH%b��%�.�������r�U�e�m�=����>�%&����ፐ�\ᮯ��S2䃝���	���d`��*�� �w�Xcr6n����I�p�#�>�,�'�tA5٪�J�9���4γ��f=c]���nz.�<�	�����	7+�nz�_��I-��-�5br5w�����+B��~~�Ưϗ 0�49c�	�Ҁ��A֣�=�s1�O��e��PQwTYY�ǔ���^�C�̹zԁ�(�3��P�~�l�'M�u>p���G{�����&�&Vn7ЃBY`c���d����2��_pqfwM˲v�%Y|#�90���{�E>�xU��9��/|�_^�(Z���Rd�[��;Yx�B�"^w�£��d~��+�X��IY���a�l��>9�}�̟�G3Rqn��	�����]$ԋ�A�����dM�@1a�5&Z�j�H���c�������]�̳�-�{4D��^��J�;�����?�Z=S>��W/Ƭ�[.�,�̵���hd��7Ó�t��OO+�=}�W���� �8rR~t�HXv�kvu�(�}�����)o��ˠv>��+�q���1LC�(�@D*� �q���(��#;��NI�ҒΟN��盪�1d=F�����G9")Ȍ���#哙M���轣��+�W-j<#��7d����k����YU3����"Tho�&W��i��4:�C���:�.P�3��0Chf��WL� ��c�HfO�Va�����fZk^E��Ư:�ZU����C܄�&͘0��Ȋ94�g�J��WJ�傲mU"c�-ǭ�8�A����<�n+���\�"̬�豊v)
/��R�_=+8` ��<,f���bn��~����)T	��P�\y&�n�V_��}�Q��� �̥�u}����%pbՋ�d*��YQ����p����mE�5^����jx���|�'��m�z��y�߸�T�H�3�S����Π�P��/ͥI�D�s���rc���w���}.����ŗ�*�c���{�J1�]����\�7�u��>G��%O�?J�$ �c�c�8�_�$������H�����;d��.�j��ŉ��A�c���LwZX�?��TBj���
m�`��660�/����I�~Q�����0]A)�#�Ki+v��޳@�!�1�����Ƀ?����te# ��%��du_Xw���N��5��Jڵ���S�
�C��Xj���p`���ռ�+�*ige1�����Y���z<?2�Z�R���¢�5t1�F�*Na
q ߔ���>l<�N� ��I�"�MiI�®�y�XN+���w�]��f�X��x<�ނ��������̄�\�����mX4�B�R��@�G]z��tCP�!���*���9���B�t�:kfǎ�!�m�݃���6{�6X7�"`��b��+����G��T�ЊgEwq�~:���(jYHC>��]��ɵ�O<g=�#Q�T<��y��e��\����#����0C��H�J��y(YoUAR4G�+��ת����X]�Ԭ!�҂w�`��G�Jo-I�STǕ�R4G1�>ك��[�3�z�k�1;zω��8>�K��k2�J�Ū�+�0�׿�'膅�i�Ɇ� d��+3�¤1S�@�v��u_�}��
��vg��.ER/�c��`{k��NB�t*���R��̾��1�H(����S?c�q&X�%e���P���ْ���'@c�ܜ�n/D�5��9b�q��W�Ml�0i��Zj9���C��Q�cA���CMT_�C'-��(ۆƙ�-�`��T��9�G܄��c@�zFi�]��;|KC6�[�����+̱M![3�3��AZ�r<�����Ϥ���sE�e=uF��3ۡ|�b��jQ\*Y�E�G<+�dM.�8&�BE-�N���;c�WP��oj٢�i��_��΄�,��%C?�\���Y��|Y�0�{��&M��ު��ӢԳW-�U�����.���N�[�����~r2���4s]I[x�������i��4GH�	z%l9@�q%�y1c� �@�r �_�4/OH��� =!Td�B&:R���l�;�12��_��su���f��M�s�S��T����9d�5JK��]W9,���/��&٭��W�L�Z��T7�Jv���_Ŵʙ��	��z���Z����FBډ�%� ]33(�`ٖ�ZW���V��G�W�!(H�$��D����[�]I�T14O�gI*o��r��}�E0w�X!����f7��.�]�c�gm�a��B�2{��8������	#Z%bv�}��;Z�z|�$Q!U[����	����/w;'����K�}�w�b�T&%RKh��]�\�[[~�)N�o�T�f�7$\��i�	z2$��q�AHP���
L����p�[D%�,�����1�ƍ�`j.Y�s(<K��gK7�- �cyBJ�x�F4���Yf��Nmy�Ą8?�1#�|���R�� >.�_���1t���I��v�s���ؙ������O�nd�w����Ǖ��]ίxy��4B�7��h	��-��������Is!�"�p���#�LS�2���@9����d�H�rpǴAIM�jc:���%+�r�Ó�v+2N��M�s��(�t��K�~���9R�7@H�9��Z��fqG!���Dw�F�ml|
�W��4ܚ��0w
�2�r�� o2�O�7�b���Ĺ��g��҄��欰�l3D���R�������U��@��C��L��,\:>,�BB\EG���.��+��2lV�~�_��'8����[���2ݑ�Dx.7�㣑%Ce�d��L���r��)���"����?N�E�h�8f�*;�2���VK�b���𣱆U�)�Пֲ����J۝���f������ϐ�?����x�7=M�?�u�T|�V?\�0\ymC%�s��5L'_%�M�����

�E
��"M����p;�H5��l�� ��S��ޯB�������]ٔ5�'��f+�U��?o��[k,�mŠ�I�U&ƾ�-�&��!��g����Ys[��v:�iS�a�7g*KK��Á�rmK����m��,�\ �|�/��<��vө�=w}}f̓�(�ܰϪ���Ӟ���%a��g��2����������&�]���N�1W]C� +��%�>Yd���UL~�+�ȝy6n��1a�R� @�b{�b��¾�nηG�=����>�^D����Ǆ6% �ѓ�L/FW��HM/ʣ)Ф=�ꀽ��;���0��b�����>��d���uߒn?_d��>�7cj��s��r0VN�����*M�Y"��=��(#��rp�?3�Cy{�6]	����>�vT�������0�0��
yѓQ�Ȥ��J�mmwp��Z�Ո�
�z�X��ڠ����p|��}�f!QƎ`���.��J7�]�l�����@X�G_
N�*���`�L&��V�S��n���E�{��3�3/��*	�W��P�9��/
����I¥�*��۟õB��݀�z~���=['�p��"��w?�&�/4'Vu�x��4�*|��Mw�9㍢��'Z�j�d1P�T ��9�뫗L	op4��+lܩ��:%�;p�n��c���a'�
�sh�����.q��9����-A�&��G�(��<��}yf�����2,c�$i-�K�Ʒu��t?�D?�ZQ,�w�nMK�W9����ԡ2����M�G�V� ��1��.�b)	����my!��5��]��܎�����<�K2�V�uk�D+&�����¸����Q�����v0W��aR��ۤ!
%������i�lИ��O���<�1g�=�xg�B���~��O�-���e9^�8����L�o��UG��[r=����� T���c�*^FS�sқ������$���-��?��;�.�%�޾�x�(�F����<�B��A�܉a���X�4!/����F���W�<�O`���ޣ�v�ԏK��͞�#�q��a���ގ[��U�vX9��M��	��z��_�`C�x�=�%�D(s���v2�u��z�Q����4���p�'"�{�$��	Jg���K�?"�Rh�v
�g��X�ƾ!�#5�&)��%�[0��^~HT�1���[��%�8�g�[o(,=�Q�'�G�*�(m�'�l#,�xk�:���S� ������GN7d8���d]P���s�2������l�k�0&��sVP��9N��Z�?H��qM.�>o}�8����&�{}2����[c?��1).fqϱ��-���<����w�W؉)�乧`�/�/��*N	;�����Z��Ҍ��y���<2}�����.�����] ��teA�l^o��_O#�n��"A��㔐�Kf���m��p_���OH�^ΐ�UJ-�5�E���֔R��H7rם�O��=��*V�Ø�J�%gr��l�O����"̮�i'/��\UN�nW��'��eE���r���*�)���ׯ�n͂{�� ��iA�@��VS.ܣr�ڟ'�=�}OT�ϊ�>�� ~�̴�B�&��P�y���Z$X:L-+�9�x3W]aZc���K�4&ke�!�:�	[�U3�xnC:�Rj0)%�:�!i�y��ˢS�ƻl~L	Ȗ:vt^B��,ën+G�еó`8�}�Ht��hѳ�G�Xⷸ��&��EYD��3z�^z���e[!�0v�pb���&��Z��>ɒ?r�h�|m;y�+�J��ZG�~J�g1^���Ѥ�ԻQےg���4�
g�l��cZ:��v�I��5��[�o�.��W�b��d�_��"�k�dk;�/��U]��y��+�G�r�r[�f,�_��W[�i�Ig)�8����$_�;��$3� V��xVu/$ɦ�f�sW�h�@����;ħՎ�-�
��7�7*�fеM	Ё����%��g*�1�KD�����j����d3-y[xc�~�cU�#�˙g���ny$ ��C����˘zm2�;�d�k �N},�Zk�$r;�����m(�}�ᭉjg��ὅ6�k��i��F���yQ����ڤ�mQuB�lJ���X�N�u���E�?6��f��	00��`���0XX�*�y�7�<Na������j�CZ�Ћ�~x�oI��&&��ű|��M�$[���ul�5���=8�k��
<�ɂ�g o��캒��������C&Exdf�Uuz圍� _\[�6ހ7H^��(�S��3�\P�!\%H�.%�*6C�U��(�-\NE�x#;�zm��a;T��:J�`[��"S��ޠ��uW�d�s`���l���2~n� �v�=Z��=ܽ:�^9*o�� }*}�[�J�+�7��Md^"���u�t]�:���Vv�x2#��&����s��Od'i^�GF�HE��P�6�'E��Հu��q�lA�O�������w�R���zW��ɻ7�7χ���k� ���I��g�xd{�W�Gr�
�������:�B2�֤ѯ_�s3�e͐�����!�N���"���
[:Ǵ=�����&;B���W��\���X�)�Xj�/�~���1Ft�jS�ً,{B��,�ě7�b�V�� +Zu,�7ɫ��ut�����v(�P&l��9�pƲ����R];� N����.��GETEN���!L6�+�Ǒ�j�����+J^hp���)רt�9u�� H�t�3O*_�g;���Qp�8�0IZ������[�f*�툉�g�L��:$*��4�/�tB�.�p �����(z�wd�WWZ{����t� F�st�lr����ݚ�%j��$vs	�W8���Ɗ��賺���}G��5<N�!��:��&�h��m��X�|<7��>��*��a�kz[�/�ŅTk ��P�Sm�9�B�X�xc��`�r�?~�_�#\q�۴xDM4�湞k�8L���E�	3{D��,-����Olt=��^����Y��r[r�J��#�,JmBC��F>�h��D����!�X�y���$$��mZ#���"��թ�u-�$��������XFκ�2�����j�?
I�^Qa�f��%Z����Q�s��%���`])7r�`F�vCOڼ�(��8��o.Y���y&���=j�}VM(�*t�a㲢�[_G*�A�P���W	�|��$Rݭ�r�U2���`g5=F|e`fp_�1�ʝ�ml�;��gJe�y.s�/;���F�l]�js�8fȑm�^��Ã�����p`d���a&��n�ӧl쭹��/�0�0��Q���J)U
��K�[Ē�(k���cY��f\r���U_l��o�+M��k�b䈥�f?�5�2�M��߻�XZt���C��i���b0��N �V%�M��DO�H�T��Z&�U^͜׵��ś�510
��,ْ���=��&��fi�/^������@��h�^���7�p#;k�h�1iq��95v�~���ބ�TFm@�F�v`14c*�9����\��#x$�Nc�h�Te�F��р��C7��4�	JQ��<W����V�۷@j���8��+ �I�F� �j���dU��I�CL��7�R���%_c���6��YP�XǾ���i��q;Z�z��C9]L;X�N*BX����}b�ڌ(I�V\6����ޖ!� ��݂�I�p������,[#i[�t?������$����UK[�m�|�wa��
8V
�U �1t�	��܈���O ����	3"�T�s�.���c�Nw�e~��u�b44�R��I3Jf��ud�cv�~: �Q|���G��y��6�aB��F�� d]\��!� ���X/�l �!���lv���
n#Q�[���q��a�V�	���,����77c]�v!n�8��W�:&Qd1B����B�q�oFH��y�$Kf�7l�u3�q�l�#d�f���X���^h�0齊P��
� ;Q�=��Pc��z��*|��r��-O��=��
�qg�*��^l���pD�H���)p�d���-�������@D��[�a����b�X ǌ8�ٛ�(��Ԣ��i�A��!��%
����so?W2j��� �3\/(Oĉ�F4t�'�2��C���xh���X�C�I2����$P��zSX����$+����"3#��W��]G7'�\|����h�<���H����u�����훆25a�B����k��3&J2ۨ���;c�/	�!U��y�)�?���o	�m�e�<:&l�;��k&�%�h2\Җ�,s�oXphە�Jd@?��&���(]nuW�'�F����K�]ӹ� �=H\�w��2�t��.�o�뀅��J���2t���ZV�z9'z���ɇ�+?�	���T�k��@�z��n�k[�v�^��}�� ���L��~�\����BK�}�?�.��
N�γ"_>�J}�*��+���q�����H�G�*B��K�s� MȞ�l��\{-"yV覆�[Ⰼ�X���'S����0�qTW#m��+i��:,�u8�O��$k�A6C��ͤ.�[�]б��^2U>t�۵�ST�l�Kr^���<����c � ӭo����et��d�٧ ��؋Y�QW��7�(�n��?�#'��d����5�İ*�9��'���8Nl5���)����RxO���0�tnz�"�G����'�e*ky�i3�Kk� NZ���T�x��5eI�׹�R�{�{J����������wt�6�|�0�CI�G¶5�0=�&`��%�ɂN�������~̏�g�z����O����I�T��C`{
7Y����J5�oA���;:���%�0;o������E��o}7�&o)S��j,A��H��⋸����|�����h���G"��õ�&�V�l3{4�z����D$���²K�o�i���?l�Uϙ�a6����ALVrX�#[w|J�)�S�iｕ�>V�" ������'�m�E��s�x���x�mӤ�svώ��*��X�KʵR�21TS��R�~�y���=*�q��"oO��۰�����z.�hnbLе2+�uU+]�J�TQ�lyrg���mE��x1߯T`�%^SY��|�E���ލtZ��l��W�j��f����_eXe2�yBt(R�q�'N\�AC�0��������QR��R���qJ�m$�p�� �%��2���j{̦��ͳf1���Xp%��.�Zۓ��q1��O?ޱt�M���c� . ���+U6�����Z��-z�Jk�@�j+�wu|b�B!�� �I�A����.Қ7��OH0S�:ԋ�,/�R|�(�c�\� =c2�Ε���ҥ����\��{�@@�L���#��ɦ�ضQdV_[f�>�T���u��P�����8#
����G����J��H�߱�__2��(�afn�:��ĠԂ�C�k�
���&R��Y<�Gcnq�{�BHG�� ��ڃ�@5O�@}肞��j�]��0��j��[g��=�m�|D�|�n �k94����D}�4rE���l���E�h�_}�N]�J&��Q
0�~3OBA�wǒ�0���7٬�︯5�q�upX���M�l�����܅�䑙YM�����ǥ������d�`1�c�^%�8Ȩ�K  �&W;4�Q�R���m�	ҺA���9Ej .����e�1�A��5�ߐ�ƕ�P�*�2�tt�X��mQU!�f��0������h�OsLbbV�^�D����@)����OC��Y��c�2�qj�6(�;�^7+ϸ���H(,�A˩�8m��1�I�@��3��O��!֛U�&V̼k��7)�D=$��|�|\�I1����m���)�$o
�V�2\nv��4�
ૢ�ѝvD`�@7�X\�rqa{q�����6y�]V+0�0/�M�7��-�سS�G����H7�'Y�eO[hNZI��m@%���\�R+������4��x�P��������O�"�XsA�_�m����]Pd:�P���$���q	�7�x�~�(%�t`R.���]�X`�w,Sϒ���P�kh;)���"F[^NY������Ű�)ڇ H��o�f󹟸�EnA���u��T��F�����.dR�-�
��3�G@�@�&E}�oŞ7�@8�����c�t�+A�,Dy���|	��r�=���SgU#�q�7�5�J�P�:��}l<�5uq��T��+��w@�s��h�(u�I�����؟�s �'� ��)�����}�}�e䧬�� ��l:9~�9�7�w�U�ֲ�w�%c��54���I,���t��6H��V1����p����9�K>�0�[���;P�s����d�-��r��jr��ӄ8^��_	;�"���M*b��=�J�HPUS����
�k ꑏ�F�L��zp�=���[ɲ��8�s@���U��;!�V�۝pW?%���}��sD��D�^^���1p���`		�6�<��gT~�9�=}('''�.y�փ5l��V�(���l*�bn�2\瓪\'�Nl�	�&����:��v�=��e�<�ν��!$��>��:��p�y{tX��P��Dat��[uf�����H�F���Ӣ6�PRk ���nn��,j��U:hg��{�VI��H���5Dg��ł��ޟ߽��*�2Kef��g����u�nu��L����$�A��V�Lӎ�rF�q��M`ԏ����3e�}�⺮�������eg��RB��:�1�b�j�����W���p�;ls�?txUD��kX��#F��T��oSw��a��||��	������@��Ic�ˣ�����,�VI�A��>��\��p�/mv�p6�~fҫ�-)�ɠ�Q/�,�1�_M����<�P"QX#�1���F*C)x��IS_�^�=ܚ"*D.O��3�fł�&U�,� �\����\��Y��M�Q3v���Al����>����&TN�u��]����͆[&-tť't�k� ��D�<bX���m��j����?���r�<�?I�7#kOZ���t�V�~��$�ŉ�5��Ӟ��uR����Qa=�b�=՛T��ǩ�"� ҽ��2�㑏|ΐ���(���쨟��Ĉ��ٱ$���i�x�ʦ����f��v�7���Ȧ:�ә�ldZ龾*fsBeo�޺	� GR��R	G_ ��Tة۰�"f/W�����v�E�JX]q~~�eq�����C�h��ϺiF���y���!ӿ͵��c���M�=����H*��^
3$���/U\I@�%���/c�`<��hҖ��F/�-�!�/���֢���M�������1y��R
r��5<Þ$iL ZM����%QGz7��>g���q��I��0���k�A���Um�_��H�TG=/���ZIb�YF"Sj��qI�q�|�Vu�Ő�ހ?s=��o���W��6&P����W��溟M��}��?�-�@�g����q�
�pjG4a��-E��'a�obV�Xca�BvU]����A�У) 4��y*�c\<fy�$�Q��>���X!�͊-�Y���������>��J���l���gH]B�0�j��@F�T%��<,v�c�Q�#W�C�S��.�cNt���`g�.KU�Ӥ^�����ɉ~#Ey	�9�[��d�$d,����T|�^���ˍ�J��eS� 9˜�����sūe�Y�7R�m��v��G��bd�|��y�c��7�Kݹc�G���5-8�������?zOm�BT6&�5	$~���߲��*̲�~��4V]9����Qk��wќ�md�mQފ�JͥZ37��N @�O���k�U������?4�:���V������zZUe�Q E��F��	I#V�V�*��-c�ř�ՙa���"=ĸ�/�>�8纐��#���)������*���8N�9X�@`��ܜ�T�%��5�zy:��T���7���?����'��~�ɣQT$/q��FW����S����b��pa�M�+!ى�vZQ�u,O][?�����/�~nk�	�ǝ�s"B�������G��~�؊_��^���<LɿJWC�M	y�O5�+2h�Pq-5o�����S������Q����13�c=�c
�Xt���n"�і��If�ݩ�0��1����������SZX7m����B:��"��Ȯ�,���m%�Id�Γ�<J��+�%�2�{t���P`�y�$;��f������zd8.C�hxY98�'�F��c	�H~�O;�W��b =���[���n"��yѭ�����	�p��'�i%�����u$p�ڜ#��/5�g�c�'��졻W�3^����`�i�o/eCV������ �d<P��%BD�>��]X�T�,��V���@#�+$#y���ٮ��9���|�Y`��ʇ�L����z3Q�s��$F�� �	�+gw"���S�ե��b����R�.��S�-h�VBEE^�(�ăT��B��B�k�|���A��
P���N�sN��K�6Jc1��ݾ@���a��Sƅ��G�i�Q'a��ղ[D2a�g�n)��ꚭ�����Yh�۷�P��G�?�
��}�^�Őp!^���N��ar�gG�#έۅP���d�=�;�߮#��D���+�Jjg�g�8�뿱�;O9?���v���U�� � ���\ 8B����u�[8�����������+�Yu�H)���d��T�0��U����{�Pm�G�h#��X��^,t�HD�mYћ��B!���u 6@�#�SU*��p>�	j���p\����]�_/�9�E�������wmLO�f�Z�<�9�e�mx�J/yu�wB��p#F���g�?>u�t��@\A,���PA8��mYѪ�9k��=�k��@�Km$�U�@��X�I�;4	�(4�:����bsf��L�YI��o�H�X��!Ը8{�(I++�x���j���m��x�}�8�ףL�2�(ދ�7�^�7A�PA�iʬs�\�K�Ȏ(lʨ��?4 �Lz����RU�-4������I`��Z������k6͌?�2���p�����Pg����Y�=W��3���/�Mνg�QZ~���'d���Eq�Y�F�\/�#8tӸ����5D�g�wvlv��ϱ�3����T"�d3��	�\��⋡���B����iumO�c�TZ������p;lX�&�Y�&h�>�rIƒ�!�3��e iy��M�J�x���S	���5�;�,�ͻN�m �c7�p sQ�ό��z�j-�������YJd�K�^����0s���Z�}�B�����o�"���lz&l8K,jrFX��ؙ#2�G�O,>.�M�k�m����P��{��e'�$�CcV�^����\Ш�Y�(���[�p�LGd�D�㏘��l����Ҕ���iط}�D%� ^�R'���h��,D�xK։\0[�q���XxF�3#��_#K���f�� W�Z�s�2ӄ��=�xB��ߨg���1'���挰��R�b�Ne�S#<�� [o��WҨ	�Yg�eV�&�ڌD�*�Z�6 ��*����>jde�g�%��Zr(dJ:f|��ђ�Ɩ�jEӶ!M�fK+%�',.� qa�1�m�Lzr��D���M�? e�/0u@T�������n)z�߷.�Uӛ���7P��d.� �}=��`a���wq��x�E�3���Ӱw�F!$�L�RI�������7w�A��w�܅���H����oFŵu4�np�_+V'#���A%�bxv����!��8�}*N�����k4�RŘ�ZR2�-���ih��q��j�@�`˼������>g=j�{�޶"wb1pHTAov��l�쟛mz� e��#�Z ��i�h��D�mU{H�7��Ip�Pa]��odxh���D�ݚg�#_Bƣ���ryed5�+�)a�MnEk-��|�D�!� ��A�#j�x�a�Z\��LS������f�N�mM"� ��T���+Y�<��u��'b��uh�A���8�E��ХT��L�Z]���c���l�&��N��9�ى����Ƒ�jk���DZҜ6-�\�� Lr Ⓦ0�([�D'�ٔ�ޱ_�2[��:�+_j����Ȗ�¢�I���J���BF� �]$��.���L8>������)G�oҝ,��7;ޟ!o��Lh���[aJ%E��
"e�Bc0��'�Oŝ?-�=},	����7�3�Q�2wj~��o���I(������u�Ўq����e�߲�/�Yu9��eC,8��~Jc�6W�5S3~N՟Q��S��υ���A�_���y���mDI��)�pC|�"97d�>V	61�j�ܪv�?(���n/"�T"�W���b����JC�"������0��@ǌ�����۲�����,��J;H�C��2N��\7S뀼�m��5(�Yt-��%{�n�H�Zo�e�k��g�����?�����:�ú�Qq���4Q�����,�Z�&�F7���(҅n㳠��L0�y�P��� &�ӵ:)r./�!!*��z�+��Y����1 �Ph��GONt�B�gx�F�l"NA�]�^�^i�?�$�핖�c�e�^������"K�@���z�@?w�c~_�e�g�>nM�8����~1M�)X^*�Go���TE���[������TK�����l��ݤ�.��mJ,n�f��-��o+YH��lSF�D<Ev�H��Ѭθ�*>�+z�~�z�:�U�bAeV�ֿ1�]*,��ҰwcP��mY#�0�r_׼KǪ->��p�	P(�$�e��)͑Bx��T�m3����%�A��+c�
�4w���������j�1{4��ָ�	6�.��A���o���ّ���� ם��u��a�o�9Os���u�
+�M�]6�Cᘁ*4�p��$p=R�]Cr�_X��+���K�Lٴ��]����E���$UA>�n*�P�{�$��0���ʪ)M>��D��h:7�� �B�9��?4�ƪt-�v%/����h_,�w`lb���su{��f@Rg��ҫv�4��3��� �W������>�u�M,����6��f�]?�\�P���xI �v.e%�H�G���a��8�:�߷�%�����<	����_�SuuZs�y۲=-Gm� I��E��^c�1�.�z�"{�|�| �ҏ'��"GUsٶ[�Ж�[Q��4ӊ��0�\�0�����Bȵ-c��24�
V�wXvAN=�:�N�"�P�Yua)pX�\h/ܳ�7�{����UG�X;�u׉P9��וg��V"���b9��~.���0��ٺ�^�EC�S�iE�-l%;X!�ܱ
�/���b?����	D���D���	��& �\l�ɕ��M�8�v�s�-j�K�n��m��xd�&x�>�Uq���C6�4��W�g�ԫ%Tk���2�ݻ�ݎ�{�g%�ǒۃ2����$A�u��s@�L�5�b�'��օ�y7���c!<�8�əC]r���z���hv��6��G�8 �,��d��Xॕ������*I�E��[`-Ḿj���р�v�?��kl�w^^cO�I��k7������3ߖ-��apzRo��T���ȂF�;�����H��@�����1)7�i=:�Z��d\=�>&O�d���8b�hܩ	�V9+��'�5(��9�F1jն���m[�ЮcE``�^B�\sc����G�� 뾅[�F�,�+O�8ؚ#���v�:�A���]�FS⵮]���i��S΁`˵ X��F��qq���������6����" ~���kUw���?��p��,00�]��9c��V�D'8S��D��t�ѿ=}>)z��C��_���v�!��({�1uL�7��k:Er�d��=>&���
4S��*A��H�n�����iq�I���x��2�3���F#�`p�Z��M�XFT[��)%Z��?�Cko��!�f�I��C��Kw4?g,�s�?�aĢ�EU=������Uٌ��T��Q��R���� cÙP��N]��ѺДp�f��5,%e�A�;R�u;P�yA�r��m�=�W2/�$���������' ��俢�Y�OQ��	֤�P�%/��CG ���n�6��HS�ʢg�JG�H�R �4�O���pb�~�;*��V�$��o[��O��^�4� y�3BQ)����*`]��S  N��~2#�$��z�bh���1��F%��wM���>q5te+`L��Ï�~7 ��⠘����RR]A"D"�������N.		N�����Ȳ��'�����g��-�a��08�V�����pdǴ��K�b �ͷa�.�q'Ei���Q���
B^�+"�a�u����
��Û8gFq����x8��mS���7�o��f���n�#��w׆�F��4r�m�:������(���Oj{IWl�2ԁE7��ȣ�ȕ�'�3!܋#};�p�:l�<6#.Q�*�us@u�&���a@>$(�9��@���w�|�Ҵs|�]+�����w
VX�|z���C�xd5���򽟮6�'�#�V͒��ka2��Trxb�!�0���|���M}k��jF��n>�?3Y%P�i=䨍%��r�R35+v�/��wrz�t��+�Jv=+�)L�Od����q<G����D�n�n���ڛ�A���[X1���&�-%�l6�蝷[�h~��0�¬H�¥�"ӄzM�>K�k�gDWW�����`�j����7U��f,J�`�-�Y�(B�T�$d0��I:2���iE�Зl�qN�q�J�/L�Ǫ��E��+�
��˸���ú�8kXk��߶��؟OSgj�!m���
��i�u����,�#od�ӟ����sgAs�o�����5	G���6c<T���^<��Sp��͗�P�t��*�H��Eӏ$Wg�]a����H�*���a�z�[A*��O�ߞ I,.�ޱTpa~��	�Il��� �����������ծ��
���0nxp�<~J�ϫ��҆��nr,�h�d����0�.�����T�����a��X��X�4�g��"(�$$w�-�I�q��|�OG����Q�m�$�ս����@�8�Pׄ��Y��I*H�2�7��r)yq�Nr7F�soe9�n;�,TE�+Ԡ��OT�q�y(��&̒]7d�n��U�<����6��]F݉� Px�$� �幒���ST���cHx��w梮}d$��ƶ]�� ��(8_�2�F��O-FY<Iv���5�4���C�̵���ϽB`��M�]��!Faj΀p��eX[�}Ihl���iV�c�L�s<��<+�9�	�.��K�q����1r��a��d���T���VOb����A���N��1����v+F	�T�(�E+�,�z�[|�y{�b��&qTD�?�!E&7P9j-��[ؙӶ㧛Bi�/:=���c,�9$Ov#��R(�k�P� Y������XG�i�Yb
�b�+��J���(i�:�!y�gQ�\�Ϋ�ŬmQ�@��(*ǹ=������W�и.C:��l��G�,NuE\�m��3,�q�;����[jV1��l��1�0�W(���v�(_;�(8.g5���8?�f#�i�U '�#U���O��F����7��E#�;Ju��z�e�s>��4Je�v��b��l�;����h0�_� ��`�J�c�~�'���6s��y��x8p,a�Y�Z��]EW���0����FG>�&�	�b9~M��4傃�x:�w��-Ѡ��@z7�r���q?Z��L��^�a���H�.T�V���2f�)�e߄Y%vI#]<F#��~&85B�",��@�H����e&�������Q��e����v�BLLf]U0�
�:Vq5��%a��9���9�����s���Z[� %J�R|uc��$ ��奮�/O�Q���*@���1��<GJT�kb~d�
ob����K���<Ci�_X�������p�mכ�'Qt�&}��g��Rr+�%�^ER^$��t?�r��<nzPd2�������:I�R�툒O��=����t�H��o7�8�B�f�s<(�O! �O힕�b{J[^�8�Lk�N��Y�"l,�[�)�����A�{�xƲN0j,g?�Y�3n�/Fc�J“����w��%B�����΋�#�8Y�?��y���k�5�p�C�	���ʿz�8&�K���]��9�T&�a�Ĕ>A�5��Wٶ2=�w]/��	����3-��FP��;�ʫ0	��:eoLFi1����#�-�q&��_Fa0S���o�1K�K��2�tv1^O�K�w���.ʹx&>8��g��+4� ����@݃EZ��s9UD.D�!i<4��7ul��*�yD�=����ݑ�4g>�e�[5ά	�,gp�6t�OR#�s�8'Z|9KղT���t}Up�#�H��V�nx����\ەk"�t��M�E�p�
R<��wߥ�6yj�Eww���J�V�_H��#6��j���٦��q�����+�ĝM\��x5������?W6���I�gE�B�ݙM�:�߼]�]���z �̊��x	�<�d��χ�C1MG�b=�#���������woF��0�N��MV��hو\;�&}x|�Pn٦Z�xVR�� �����]�~�!U��Ю�j�L&��nb=w|�0@C�N�s��)0�[@Y-!J��5F��5�%0�9��8�e=�).�"�X��ܓ�{�.��${",q�)5򟤏j��ݩ�ǄXl�r5ŅhKu��H�3ԗхw,~��Q|�*��l�t���*�Aa|�3ggXX�,���W�W}$�U��2�Ƃ�h�{�KM����-K%ܛܵX,z9�kL�>]�
��ge ��*F�]�V�z0,�ީW;8��}v٠��`G�{����,�P��:�8 A%�1�cVl��G���v�(~r��f4qF�  ��q<��{�zr��2ZѭX��*��H��q��$q�R�7�I�5\�@�����ғ�1�L	�&��N�FV��ۀ�9���S��W)Ӆڢ`��A5D�[Z[���TXuY�]��S�Ǧ�X��R��߯�w�Ae%��X~����3����y��s��\}��_��y(���T�7��-qn<�1\���+w�5�TEC�K��M�R�\��E����[]��w�'����	6o,�1�dљ[C����b�<u���ԏTy^JE���AXz��n��,�rd�o6Ȫ3�!� �k��p� }��-�(���gJh��7�U��A��x�%���Y3�lt��uE�ix��/(�����9U�<Kfdi����)�`�s"�t��V5�r���;X�~�����wR���^�;_��ſ��Ӯ0�@�1H�Tx
�{#��'C�ID�α�Uߺ[i��|="WW�ِ�����if6�#���.�v�Y[�;������P�A�P4�swՓ���mx�s��Mk���!:է)x�� ���(;ڴ��LğN�K�/r(7$'�5��,T^f���ˢ�h���
��ZLГ��&=.*� j��q��,�?� 奀�k[�W9�&kS��t�L[jL+�hTB&��jǏ�]�6�@s���6��WQ��!���AZvO�V���pL��3�bJe���`�#"� c�?>��@-4g�-�־\�|]�4�z����` ��FJxu��'?۔\�_��#����� �1˿(��/9���Ϙ�6Ρ<F�r]�Zi� ���ݓPw��W���B"��)�o�ٲl�F.��>���o���&���kS&d���Xs#w�i U�|���8v��1����*��g����%��u��$�'�4)F�-}#�3�o����F����q~�р�������ޥO��o�C�d�}�Y�w7z wC�z������tct<�6�umD-Ƣu��܊�Q�z�AL�N�}lƄO1P�5\,.fF�S�8Z�"jB�
�ϜS0�$������f�\#����K��c%����خf&m��Q%w���'�~�uT����n��h�|�q爵3�P"������>�qsHݡ?�'|a�h7��]x����Z���Ŵ�W�F���I�� ��"5��oĠ*�ۀLpl��*2(�_(;�I��΄�k�"�����Ж�63
�'o_<��ܤX'7�hQ�w�!{|v�A�Α�����G�{�B����*͵�`*�*%h�tQp �c ۉͶlu_���G>��P��ચ�Wj���(��E�� �	�$�~�螻y�l6���R��ގ�?c��y��d�ha��:�<;
?ynl|�&�A�<RY�N���H��u��uV�td���Pn�]�[7S�żDLPg������#��h�c�
�6�8�A�O99�'(���3���^hu���_Q~��/r��|����C��g+n� �P�600�}s�,_Ia�EXS�^%-�j S�7�	9!�՟ l֪
�w(~�s��ϒ�����U�=o:>h"�<}�7]\��N���e��c�We��+�D?X�,��&j�r�KP\���۟R+������"8Z��e��_���Dx�pC�;����Q[��SA�v�)/�m#Q4�,A��Gg�7#��
I(R�;�.��0,��	�&Բ��/������p�<?Q��%�c�+F�01�n�'�O��
���m�e�x��5�4��F�`Ua�}����C�V�?B���b��e�f�U��̗�ec"b+\��q�ųg�*r'�Ͻ!��!��
D�!���<��I�%�8��(��Bn��#��Q�>��T��|�x�*�-Wd����f���9�p���(Jϐ�����187M��z�Q�\�6��-��z4H�'�6�@t�4�<��y�߶�*���;�v��N��MVo���hz���<���8�ԝ��@N+�H�d�����!����A �x��׌���pWf�qNS�H9�L��:���.���m�S��#l��J�	%��5��v.Օc�z���v<"�*���`���i.B c᧙��x�(vP y�Ky�s �7�<������w������%Њ#u����T0����-�ģ_ K�yf����y�\�xs��;}��Hz[Q�M|���[h��RǬ�ǾN%L����u�c(��Ju�I��t�ap[N#c�a���(��_��fۆO��h����P�;TS��t����`�Qt��������!ѧ;[��u�#�����A|c)�M[x����z�+������9���	���vo��>�e�>tS�ve��@��t���9Aۡה
H:�=��(�30~h�>�ۂ��R1���O?+�8}p=�2a��e�=a�=>uw��X!�����$��i#t��E���H�n�B��e����u�Y���&-D�C���AUn�B�~�-Q��?O�(�Y�����j~i���ϸ��J�V�Ĉ�}����*�b�=0.��{Ţ�C"hǂ�~y95rh-4F̾�mȑq�Cj���ub]�=D���y=����?-.��wIi� n��/F���٥��Skf53F�w�����G�T��!RP"��ʵ��&�WL��p��6�%���Z�M��I��ĳ-TK;1�L����jn9⏊\d�)1��%�W�	�YM4~2V���[�U��D��{�}�nc3l�Zf �R���7��%>��i"�(4��x{�p��(��y��l��ĉ������6أP��5Igt�!�Y�"���f�b�����_��ɭ���JQ�뱙h��~sa�L5��NoWj���l�L��,Ge�k(�0�Z�����M]��:9e6Y���]lot�T9$�r�]�S��<POBw!o����	��[}5`�6�B���jg,]��"��SU}D:d��\�q��Sh�����9A�����ץ�����8��x�O��bS��"����M�~Sy�P���e�~cC���a,���
*J���fe��w=�!��+b���e�3q)(쨡�!�����d��U�ƻ��+�X�3s׀9a��ܑ�v��@��:�kL�vgN���ǩz������*7Ň�/dś7FlQh�_��0�F�+^�j�����r��Pz@�˺��1�V�ji*��Ѵӝ�-3n�fX�#��:q=?�:���	y�V�~[���W�h�N7,7!t�5��Q��ڽ�����Ч�Ro����z7Ư�ǥq�-)m�|�?��S@"t���|r���I	���v�R@N^��*�>7H9!0�_$�'�D�ɪ������oO�S����.M�u��d��[X���@L)�����v�C	���%�,�a�o��8��y�|�$�ggk'��'�w���A���gX��3����zm�.�r���7"N�&O&�$�l)���`����,�B�.�%�"��}{�ԣr��@{�l|�+���	D��b����xw$�T�/;!��lF� �0�R)��v��SW��8
%�5���z{=(+[��Qn���sn���Υ=�k���T���h�h�1� g����`/�W��wa2�`�W~�{�J��=�t(cMQ��F:�;��
i����@���W�}_�Z�B�6���J�R�#�kD�
m/^��"q|e�ë1ǹ W����B���fE��g�<Q�ny�F���o�J<d�gXu�,��y��ᔻ/*�-��Yp�,k���]}_�ϝ��0�aG�v�56-���41�3ɀD>��g��ЦF'�߉>;Z�=���,v�Ɵxr��5Emj��^��=Ȋ�Ԃ�����y�v�?�o�Q7Vf��'��b`'��=�>�Դ�v�U٭��9�6���xg�8�	�����9�~�dFviXP������D~+g�O0y��՚L��������0:Dx ̹�M)o��{<H��nl�)1����fl�̵ǌ�R=����K��P�i2b�˾(;�6����ֿj'��g��b}2A�m��-��yľa}�uA	�(}b՝^o:FP�����g�Tkޏ�����h�qF3��x�b���Ow�{RPIp��K�� 
YP�Bu��j�~��Ϩ����$I��r'>���q��z$Ôk����x�#Va)v|x� $61 ����va��xLU6��!#20R�ʿ�s
�������V"��l?wݙw;�`�T.o��k�rB�y�l��J��y��8b���$��R�E�YwEhրx��ۏg��mp5l�U����ԡJ���}�����c���ҙ�=�MP�45}��� bĩ�C�����m �14 ��*��\�D��@;�O���0��`{{`��Q�4(���)�1f'x��d��i�r�w�6[��ȀRP\Ew;O�m��B�͎0��"�⅓�@�V��}��#�L겖[�ȕ+���"Kt��мߟ����y��3���@��p�4$�4�� ��%�:��4�p�-_�n��
g6��yce6VB�6�:�R=�B�)<z��&��u5�H\���>�̽��o65��f)~<лs
�P�����j��pJO�'�\bĦIK��c~>��J�R`[d�:)q��P��a��+Rh�1�-p��>����.�gND5W���O��m�E<��qc�F���Ω܃�Q��r}�P	�z�Aj^������&"u~Ƴ�7�6?�U�E:B��P���j����\^L��G�J��q|o���Br,!��лpj�ϜK�#��*/$�H$��S)�U:�̵�\PiN;�c�����\�:�����R(};���t�:�!H�V���G2���+34;$c�f�t�ޮ�
����&�}���C/�E?�����
9 eH�ɣ�Ek���||z<y.�7:� ��E]{?3hx��^:{T�Fla��X�*���r�Ꮍm)�����i/�A���ȇ�Z�3pQ� )�=�o6�]�u���(mH�g�x;#Į�`��-�1�y=��S��t���D�IWX��E��$�%>�W�X&Y��(~`����/��P.�3s.��+�l����.P	T�[J*
������,�a;_�w��&<�?�-2����]�+��Ū7���Ĕ����6F��4�.�I��c�mo����
pE/O�i��m1�=
��.c�?��ǰ~���~h����u��'�,���p�42���kYb"��u���Xwj��-�ƥ%Vu+��������_^J� �/K�s��a�Җ"�/�Q�\��#Z�����YX�7����������r5	24$�/��E&A-��C#�=?j�|*~�_�.	�d�N�osE�s>���L<p;ɪ���ݎA�]��6�@���Gl=�$̸��"�/�-�{~��8���[6��H��8L��R�}���Ws��т%&�<����uR߽��
`���qi[����ke��;��X񜽜Z�X.��Ėݫ�мQ��84M�I?6��dˮB�0����Eb��X,D"��� ��[oڜ:�F���E���&�9>	x4
^ߒ��kK'��)Q�ݶ2>q�O����⨺x.���c<B8��
}~���j��1ב��.vI|��[�ˉR��*>v�u7��O�o�3����g!-�@ @9���y�������>h?Pr@�v�F4����t�I��`�3}��L&W\x�[<�j���g�o��"�)���K�H����BA!��=?Eh���оx'͸��|b�֤ʮI�v�nk�����6[���l��1��P�F����e<�K��z�o�*�շ��M��XF32�� �� y�n�5�2�F�#�VT*ܥ���NWt��0��ҽ3MNX��Gzq��.hM�%w�i����E؝E���%��:  P�@l�-���ι�L���x�ėS�3�k{ssL�/�q��~))�R�/��w"�_��xhG�3�{��yX\Ȏ:yI]�yx�x6�qd(�;%C�Z-|����W<��/�~p2�3�N �0�N���K�Д�5)f%�Ӻc�pmwY�N�L.�3J���ڗ0��o�/� n�\�F�d�	�y$�;5+�G>�on��	I�o|<�E_!�H�++�B<Y�]sk�a��	�Gճ�3���Y=^���)�c�:��[e���cq�+Gf�@���b���c�R�I���UK������'�����o�����9`�D�����t�Ͽ�S�����is�����)#t[2��rY<��Ű-�q�kV(�@�J�al|)J2�*��^���:����*��>7�Iw��0|�z����ul� ���L'����5�J|	@%Z�?��@7�싨.����?���1��0���ՙILγ��F������ۉ�n�j��'���7~Þv�p�}e,���r�S��W� �k�� r��·�`�s�h�L+]?9��$� �E}��8�ᒶ�?�Y&v���)S#�Jg�>�Z���}Y\�4{��Z��g#'����ށ��Z�}��)���B�v�$Ry�̴j����B~��A7��u-Ƒ�d�#Z�{8��BiWƦ	RG�u�Y���c�(W�!�szF����o�Q�����!l{�d��1�k<�¬J3n36kS8I��M0�"s����2��k�Ȇ���R �
�P�|�f�je �,?+�������f�|�����|<��@	�P�����ll��|Ym��� ��z�"����� ���EdQ���`^c�Y�17�jͱ�z'�I"�̣��r6�����b�Y� S�R��7�=�\��	��(�kƴ���:�0��.��u$����4W�Q������ʋj˻0*�v��+8�O2�}S�mʜ�]敲�U�\2$��ꋕ����Z�!]]���!��.�����m���Qd �Vw��{�ӷ� 6n�����3��q�>�k�A��Kx$����%:ĥcm�sS�&��w���I����]������v����lq�{NC$�l��U>t�y3|6�
|�\\��4'�m���C���6�a}cH_ʸ�U�z�7���U�|���F����+tv�?�`��N*����3��eE\j�{E'�q=���@M6j�)�t�gǝoK���p�R:�6���W��`I��f	)X���N1|70#O p|����̋1�կX��1���r�Z����Tzk fe� ׉���s'<�Y*5�R)u:�4��ڏ�Ig�*8�AC�暸��Lm�FX$}��H,����G��bh��^�4�d��&���:d�{X��ڙ�G�-(l�H���3A���I@.&��|I� ��G]V��{V���;�q���4�����l���a��%Q��e˺K�
(L��:S������^pUE{3���(3����I��G�Q�� �ѭ{�(�{ntmM�93l��2=]�U��@>�N��o��Ka��ғUm+r#�\��+�k �N�ae��Ȍ��DT� v�g!ٔ�s��9�۝�br��<ڗ>2�����N�}�q=K<vB�s$�C���͵7�o�Z�U�mx~�~��8~�F=̌Y�aF2����x���X�9��f2\�,��F>���ïӜ�zKpU���7�/c4��T���s�렗J�+�$�ٶS JzHv�)$6(�F2L�v��Y���Q߿��.��뚧}C�%N	c3�����a�W�~��ſ�Q���W��Q�1fx�����Q?���4�5u;��?�=Ȥ�{�c���jG3��;[���z�̹.�r�-�غ=I�����gf(�G�w�?���z��leZ�U��͡�M~9��+>�|�E@]J+��x�O����>����}�Z�53%\�-#y^�Z�e1ķ�~�oO4���?����g��5�0�Rl��Ϋ9nJƯ?|{�����ӒC�jJEt�����J�Y���4�_)��%��a�G��$Fͨ!�Y�N�M�l��J���9-�� �5��8�����CZ���ʗV��3����Y��`ӽ�||�kZ��䥾�pϋو˞t����4rK�+%��2�3�ȴ=�³0sQ ���le~>��)�O(n��l���'������>�A�V�.9Fz��w[�h��{��AA�%�L~�[��}���l��>ow�<�YC��B�03����c��߮��,|�$��][����c�I�~�U��Xz�uzĦ��������C)�(�Ō��.	�ڧ[tOF�^Q��"Bn0cy5m�Ӥ]�[	�;:SX�0����^z>��N���""�߮jU��ͧ�j��}���6�z=����Zi�ia�-��;�Y���4!�]C٭L�zIj0�o5���L����&�����l���ԡ�E���WY��� �;؀SWR "�mVxtG_�@M67mK0�(�w����#���m�NQDZ2�_�yխ����6���:+���Yu�$� %��@w�sg/��Xy{K�?�r'L��Q��f�v�s�Ǥ��KE?���*_<~�>1�u#-���1.7���Ru��ـ�[��[��y�:M'��Y;H�2�r檕����}k%�t�;������a��C�Ih�pߛ��R��P����6NR��-[����[��1��~�v���<�6� :��:��&�C��DIC3�!�;Z�+�|*p�|���EH3l�XBZ�1��d�J�j6چ�Ss�~v��>���|h�W�I��YϏ(��^�ړ�(S�Ö���_�ly��&�D��Y���m�HK&C�rF1�(��5C����z+{a��Ld�s�=�g1/W2=��Gk�5Z�an���t{������D�*��~x�lrq��*�
�RP4����\��bQ49޺�ÆifE:O�K�.]E2�+;�nm_� |�Β}x˦��轡�
�C'B��յ�� �u^GF�^����oT�hDь}��@Ý@)��R�3�>�c�}� 6,,,���
>gIZ��Ve$#���0�(�c��ɼ˩��LW�+�r�h��
v����j���d�z�Xt<`�:��%;v4���	��	�WrA���%�o������ldk�yh��9��0��!���<P��`� {T������1��]H���Bog)<Ks���0��_�����fG�rߵ�Z�7�ոZ��	�Q��'/g��'�f0��%�]hB˫�
1�?�!Md4������K7��ݾ��od����E�u�������툰���o�܁ �����@o.��Ŝ�Y4<�Ֆ{�#3k���lG�� �!��L��Ǭݿ���jF�����+E��PPJdʿ��HM!=�aE<9ӑ�o�@`R���WSw�t��c���9�V	�>�v�<�9XU�<����-D�u&m,pԏ���MnK3|���pV�6ws�����C�k15WR4p5�Q)���'�*��/:���dFjTC[V����=ua
$���T ����D_G��PMc��'Hp#Cb�hE�	�i����òf�>_�A'���ț���<'��~�Z'!\[s/'n_N��#0�x[2��^.����Z�"��X�A��[�c�(+Dqk���g��!�7b���g@�������hHaw�����m�2vf,�ERJ]�s���@�T�MB(�FYu]-����ydDM����v���h1��GF2��'I#F4;y�5_�h��NR�N�`��E�R?��ղ�ww��0��]q�h��¡X�^7�~�4�aV�]�<�]I�ry���'~/���#ޗJ(�-\l��u�ߥ��l��h����g�[�T��p��wD��WT�x���7ٽ/�Ŕ�jP�"u�ɉ7�*��a.���8�Հ̠:!u�c;��P>���\T���n"�<	�è:4\9���e\�����=��gP��m-�yCC�hY*�8�9[I#��F�N
�����ԛ�6�z�7_<2��c�ʍ��Q̭�.n�6b|w��gC��*�v�����(}z���jV0Ѻ����s��l�"j�o�upt�����i0UHn�F���{Tg�<����Āj�ew���2o�M>G��X���!��1We��°b��oJO���H'@?Gސ�̭ަkb֙��H���B����x�2�r���H�$<&�+^��UR�6����ǹ�*�����UW��߇@A`R�s����rFp�*������Q[X�;�o�Kt�pQlI���:e߷Y��� �Z�Ͼ�6�,����syS�O������D�}"�Ac��o���S
��@�}�t`E,�z��e �l�)yf��Y@X@(�4�$ڛ��L��6�H��=9�hY9��6U��@�"��{���3��?9j*D2�yY� ko�.t�v�'��AF�� �ܰ[�I�1�0z� ���F����I�[�"�l�!�;�H/�[�b�3�����O;�{ѫ_ThQD-	G+A虼X�#x,4�i������Z��{�S0{ &���d�r���[l�,�p��R{����ʊ���^��ݼ�@��^��(�h�=�F��F�.y��a��
/�n���n�Q*��J6]Y�5J���K]h�sM��B����W(%��S�V�<�Q3�1���;ݕ;HT� ��z�*Xupx� ��#?Ҿ��*p-�j��o��F8��06��vp�х�l�ɱ���|��ơ`, lu��B2�����h��nc0d��i9�����|��rdZ�K0 �O�[R@8rt-���ަ�g��A�#Z��ω1kq�ȸ� ��r�ޚ�d�+�� �N}Pll�s��y��7xi��bn8�m��2���J1J_���Ŀ��3�F<��"_L:�%ʎ�Y^�7�2�������8���"�-��l�	�M�S��<	?R�/o��T����ɸ)��7]I.n\tu�4���n	~���4yyc��9�׉��ٜ�;R�!ѩ��,�Ca�wYK��ِ')C�eZ��٧6���̺3'f��8�!ϧS�$�I�{�y�7>�&��1�_6�Ư��	 �y��Ш�;4��'X$�����o/��E�e�J��/I\I�i+�S��[R���r"S����F�~��\M?��K��l%�
c����k,�G�o����xnnT6(�+wՔ%�	_<�>���;������M&��P�Ko-.xW s
^��[�އ�NH]
U���9]$��b�Nj��i���Xs�I���0�5O���r�r�і�и�F��Y�]u���RC���U����1�<��E�%(<x�[�2�̭_F�xH^5�o;�ɜ,�9�/���;�yyY�_���a���$�SC�+�}�����aV]H�ږKЉgN	i���h�Y���[	����z2�%j�Y�{��<Mt����X���:��,���)�x���h{!�O�~����O��t��o��@=|���)�
��Lt�G�fK��Z9(J�V}`���_:Iy9}�^Z�%�0�����5K�����I��v�H�PQ�jiN�=�A��㒘F�ZٿN)� H��) ���@�D�)"�\�>�������EET�I�Q�6��W�����@��4�dq�74Ѽ���.G�t�*\A
�?}�e}A������E�L�}�0#�t��R�Q�z��G�K�,���)Ԇ=۩�8�U��ث��(�V��IH�-gf���W����X9�ɢ�a���\ā���1�c/��r�]S\ń��>F|�rDl�7GI�ۥۋL�����$v�d������Ptm����Ɩ�2A~�h��S5JvHCɋ'���89����y!L�e��j�Q۶�����e^̯��p,�k{�����>���\W�Q��~("����L'^�Td�jb�Mn����ۻ�D�����7L_�;��d-h+��~�MHE�n�U8�e�Eq)��-�r3��ۼ6:ܠ֕T�o>��2�da3����O'0vno�S>���p8�Y�Uj2f�i�L=2a|=Y&�$[�P�R�R4����W�Y�}�+c���z����Q���E�לm8kŇui�f1)6��(�x���c-�TkS{�gьN�����?�G$g-�p��ڒ��2��&�,.�cF��i�|}�d0�zP��m�4�H�k~�ӻ\9��3����֨���&T�\My[���2'����v�ī	���=��.�땡MX���0S�'A'�+b��}B�V�eUv�۲�7v��=QDg�g^���bdP��	��?։�@�6���h�LX�@V����]`nȟc�mв�}���_�h����x���foS�v�o��U[��F*�\9u����AyY�6'���u:B��/����i�5,��'�!>؋��&� X�����Ϩg1>|}���DY�1�ܒ~�Vc�u�c	�#Q�5B�o�}ܾ����p��+,4$���j~**~s�I�ݝ,��R�L$��A�Z=�e��D��3/X�~G�o�Q�/���[�v_�;S��9�8ա�NS�m%oX/|��z�Xl��!��K�D[QB��$Q8q�'�o�נ��V߽c��{�_�r������G�_Q=Qݭ�1��D�==�LJV�ǉ�������_�ko��H�m=����-�q1�< �4��uHoiU+��m�c�/yB�N
�RB�hU�kk�L�qy�X�6̧tEQ�ϭ�bl��>�\�T��6(�42x���S}r���ʖ,'�
�W"7�k�]��ӭ�um-�8�|��b�ݟ^4i�Ho�Rn\�����)�E�x�h{���O�6?�J ��ɇX<)=���|K������n����e���ۂ�xW6����=<���h���Ue%�p���;oC��*������ex�8.�"�^5I��ͤ�tm�i1�+��*�Q�<(��<|�@M�re���,enxR/)�T=k��[�U�e1�_
�~�8 ?�:p�H������܉We�����:��*1��f�5=Q���ڛ���G�H�ٔIڭ[ nl�;���\^�s���Ǣ
���Vw	��dMMY.�����xTc�^�q-oJ� �c���J�*˦aWH��z�b�����p�d�U�7�
�������u�|R��c�)^7�3bXD9�V�8�.�p��f��LO;-1�"o���eC��?{t2�$\D\D�2ᑞA5���6Ǥ+_��o?�4| ϼoz��������GH L�jB�vk5��6r�ӈ��f�N����Y4��ŕ�e�Ve�x�j9X�s�Qҭ�i(_��&2:�Z�	��? 6��f���\W�maJ)M,[4�2���7=���"&D+��b�!@l*��{%�6� su��p�~J#%������>�2F��ˀcn�H.��_@�Dg<T��a庂��.�cnK�<��2j��ʭ����V।Z���)���D"��t	�l�<�1&�-���S�G�b(�"\P��1`<O�����!~z�_�kO���g铔��y��tz6%��ߣ>�@@����%�S�y=8a�Tx�����3��"	"H1���+v��4�ZW�(#="��g+�o����g��AF���OX������ J�	|y�~����x�*�����'Оڸ�!�~xc����K��7sv�X�`4���+��y9�8��xg3�/����A�7y_`�����T^��7V�׋!8I�N@��)~ħ,/���G"��E��eS��L��cz��!n`T3�!��L�NX��L:�F)��g	q+�s�g��q���X��ёതE�ZuS��,�	���S��T��X�u�ͽ���!�R,�����>�A7�u:c���q��X�g=V�=rui�X��AJ˓�FȤb��O�sN�o��,�����B.�?s]į�ǩ+���8�3��3x3_3[��k�N����n퇍d�D�Ow��1�����w2��6fU�ub0ٔa���<e&בkτIZ�v��udw0��i5�;��\go���k �R�҇h]��,6��aXЧ���Zm؍`�k���Cܤ��6S	c���n�~�n�|k�B�	n�����P	��i~f�Nfq繉kT��K���\���і$���a���F!�։��� nEN{������'�V��A?�<�!��G@�v����aS�y1��=��R��gs�L��і� ��u�2������#[	3j��k7��x���:���4�o�!�QNM�ڣӣ���<�.(��6�6�a������p����{GAjj�	�8� n� Rߐ��P0x��/�hڌ����u[E^���|�`V��,[�64�k��r7���*M!v����Ε>i��`�[w	����S\��%�*ڛu�4�9���]�j���Am0[���C_�RM�/	�0u��Qo�Ӟ����������T�ɯ�Od�c�@>s]��+�>"_0?�+��z`������"�����:�\����Rz�#3��,��b��=�	��A��}��/"���IⒼY��Ԝ�(�;����"�{�n}�B�&��b�7�\;��R���	~&�)qM������I��X�9���h��Sն�HE�����(ݳ��`5�NJ�(�s�sy�I�6��6岮VQx�D!��"�c���,� x�"~����:n����o\�|E����#�L��_�&Fm���'��/�޻Ԛ�D-�d��#�U���U������͉g�&-�d��<\���
�-e\����T<V�:2����з�3�ߛ����E4w~�{�{,%��ڌɱ��D�[e�y�5�X�`%R���<��W9��B���]�ےnO�fȐ*����#�U>�#Lh��@�[Xl�.M9�ǻ.!KS,�L��,Qw���	�1���b3ˢ���'��Tl[�����v���"�~���HÐ��*κ�Vc\�����FBG��7@�i�RM� k5��/�a�d/���Q���&�-�W��U��/��-0T�:ȶ�����֊�c�U������-��X��Z��~�;	����E���Z��Ԓ�eX1�_t�i��� ����,���ϝ��;�x�[)�9E,9���V��9���� ���"~ph����F��<κa�C�
�M�%�b�_K����%�Xk���-/��8�;�����uRِ�	��x<Ʌ��#��;h]}Yy��|��s�0!�����gFy�9,B�*�]g���V�g}1���@�:�I#�?\�(�ϗhP�l)�����Da�
.��I���]�Ge2;MI�����N@����+A5o=�j�3�4�+-��5 g@�����u�Ӧ��g�,&?8{s_ æ1k6�
UU�W}40�J8��.���UM��NSewC���k��,���F�u�n�ֿj����* -/���pS^LD�)%���@(�Ч�f��SI���aߑ�5��F��$a�W��K�YN�����F�K��C���*�Q���/�󞙎��.�d�^���>�+c�(E�䋴k�[�?��Ӆ��S`�q!\� [���"g�9�v�Y�7�`s]7�#T����%�V2ڗ7b�(8��N���<*�.y�́K���k�5�S>����Z$L��0�Uy�*Wu���S��ګv�Ӌ��m9�;�v��b�:��12��|��^MK�d3��M}Q���ZLV*�iH�eH�B�R`)��wLc���hl��F���4Nw$�l����q+�0T^��S�E�G�5�����N���^;�p?��M�_P�
����Y�=C�V�-��X�q$����3�S�F�J��7�ዩ'���.�e�=|�Kx��?���T�����>a[F�XR%v����������z3�=�5d�s*u����Au���c2?k��<-����^�E�P"3�Cƹ�
ߣ̽�H}%�.�(�{{����/BȌl#�M̎���:�>@Or'��!��|����k�$�qҫ�j�����AH`�61�_�j�F�������j@���]^<�ɴ�L�.�xj<Q��X��`�m�~e+��y�F�y[[[ B2J��]d�����f4�p�^�k�G�i�Tm�mS�PtSP�"e�)F�b�)n��-�j׃��C�:s �aY�U=eg���1���=>D����������IN��y�y!�.(L��엯|w��X�2�~n�}��ҽ.)�Y],�΢T�h����^����&������ջ�l�#t��!<s���@Ut"nأ>�.��;0ÃC�%�!)1�C�vC�}���r��90����ϟ��M�n�ՠE�C��,��T���v�O^�x(��1$C��R?D��j�S����rƹ�r��	3]ZX�>��E]�
p`L<_w�J.��q9��[J�	�iT����C�&����l(Px��Pܬ�Q������+8`�Prs��9���a&�j2�>� \�<OvB��2ttl�7�&�Z��R��!���]V�l�Ր)-遲����Y@H�|S;�{^j)���.�t��$�q|!�?v_�K�w�VM�Z����,��2�W|navJ*g�H�P��4�o�U�S��7���'����l�׭�1A�W�m�B�g���1�1�bR�y�׮�_�`R�EI���I��] �]K:�� �6˯����D`H?���`jil~�!�_&n�\Iy!�!%#l�YOF'6�x_��#)t��2�Cv�$�i*B6Ⱥ�4�'ŭAQ�G�����2�~���.�<����-�4���8���Y]�N<��c0D��*���宨��v��]\��"��`F�]�?ˈu��/'�}ے.�(BE���|E�)��+t[<Vܳ?�rPJ:R_^ٛ����r��|�G:'�ٓ�� x��J W���.P^8��~k������Taq��c�T�j�� �%��?AģA-*�*B(�W+�LI<��T��VhHP��:�Z�˴�m��A��c�0Hlj������^p��P1���� ���O�Qh�Is���Hlnf�f6�<�2�]�H�M�W�q\�ˮ�\�4Bwײ��h��L�����7���e��!ξJ#�$Z����tb�'n|й</��{�K� sa䐧^�Ϥ�|5�A�A�l߇Fjd��%�ȳ��{H8F���[�
�#p߿c�^w�>�{n�\��$ژ	-`yc&nx�d�dt��Up�����đ�91��^�}T�c���"��1���%)��`�qg
(*j�	f���Τ� \;�j���L�� ��<�~؄�j3�'�R-��25��i7�suM3ZN�9�d�$q�\�����xH?]p��03�# ��Cdr�zA��wV1S
q`��#t�p��[�������O��w�ӌе�(�<o��2��lO�7M(��^���|�n*&��ԫt$Q$Q��nKόw�e�;�ԡ�ԩ��5krz�Ч�}�䰚F�U�:Ҭ�A��۾`���f I�1N������#�S*{Qb=$G�y�Z��8�,��a��L�Һ��B�"�R�ƽM�����O-�(� �m��x�۬�,����	����>��%�@�׌!�y#�E�5*�z"ӫf�����7֓ܮ
��,�L?��l��i�[�C٪�wp�<?�{|�C�;(�VZoM�J��p�ܠU2���t�Ĵ[�@ Ln2$O]�W�AN+�Y�@'Ӕ��B1�O~�!��������%c�FE�b�[����D̶��9>e�'��� �|7o���;�@B��M]@�Z� ��Ǥ�����ږ2Y�Kg����b5g��M�&7'��񠩇ic�3�*�KU��
����O�L�/�94�%����A�t���4��o��B1��7��^V�l�'��2�S��P8~<���O����2���4���%�jiZ��W�/}KC6,�.��"Y�rB@Z<$m�51LEkHI'`@�)��B�D��j��\�J�x6q�rO��*	����Gnn����[b��i�o�}�8�0z��\� L�Z2��)��2�r~"5G�LEJ�fd�6b�D��P�2.&�&u��`����q%��p�dcs��p*��r�󯭤7�����uCm� �g�=3�]�7B�˗Q��[.z�����O6�D��\��rkG�"�֣:J�ˉ͇g�+���f��/m��Pmfޑ��ɑ��H�ꁩ�ʋ�Nħ�)T٢�l�)��PU���)�Ƣn�w��̼���W��c鑽��a�M��B��'�.A�K�{�ߤ�W������ot	M��H8�/�g��ѷ�"�85����F�G��R��<F0i���.iֺ=�U�����E�����]�^<nɗ?}�4mbm��-� ������ v�XO��m��yu��ke/���+��b�@���/iH:���_���sp%�$ ��e�N�ñާX����I��*�d�'�b;"�����_���>TW`�U��| ����%���YS�H.�'��%I�Do�ԟ��w�����m�M�Hҁ���f���0I^�d$Zf��.��cJ�@t�"��}�*V_D��k˚�<�0�X�����0�e�X��1��f����b_-��\ѱ? VHY�R�)����� �2�U��M�x��&8�ŁoR��w��\���ٿ�v�w۷=)�ƼB���(�9��:�cМ5��Ա )�ܗ\/��~�A��<���u22�m��ڨ?Aa~��2B����~`��K�f`��+�E��~s6�֌h�f�7V�8���$#���	W*W
��/��٫Y���9���{�-V�0���K��J��A�ZM��\~���]���j� =���ŀA���o�M�8f��\Y��I�ʵ�B"��f��Gm��;d��2��|^#:p�%���d���������~�&��8d�CM�^�T�O���M_�ī7ׇ�M����/ē���`�'yO����Y��1�T�V^v��i�˹�F"�|A͇�юw�+6���C�P=�Jg�{�r�=��pǕ�R\�)��U@�<�xa�ƏV�W��av˿��k|�m�a�gMmMj�BKBY�~�3�b�pu|&�����J�"��Ý(.Y�iA�|YhH�C���1|X��*]����b��P���q/$�s�Qq��V�����S
8p��q萻c��gf(�Ot�4�[�-�n�ڲ�0#�̒�n*!���WUpD���S=�-؟烚=�2����F����Q&�6V�b6p��1���P�vY%�gE�/ho.��?L*�9!�B�tP���6��ᰲ��){�s������"�W��D^w.;�2�J�h��z���>r����X�6#�2?����ށ/%�#��9J���AIi��n8�_W�����K��$�\���a �7�Ӏ�tl�(�5	�56���{F(3��rT�}4���t1�ɔ��J��{����G޴.��b9DG���zu���|�j �4X@��ʬ��;X�y�z��Y��~JKC�S�ca��5�>Oĥ�L���>t�kqo�	)/ri�`��h�[q��Oշ�������ᆰm�Vyɉ��e��<(5c��X;<Ԛ\������im�x|����sn��E0���m���39 �Ky'��aI?�(��Gϲ�I]Sa��f���u�5W�Lڬ���SbQ	3�!\iGJ%lO�)��h̘��,�9O�)ܝj�dɒ��UG5g�����Ooם�@��SE�3S��z����L���Åλ�=}�<HFu����Ek���o�A����b��`(����O��J-h��z��CD,$�,|{����H�6�^�����:5b5���v���]�0 ߎ�ۭU�P+9���ˈ���R`�8�s��3l�Ϋ�[U��(9t�̓��"�:e���c|Ti�&��:x0?����W���n��#L&�u������gű�b4���6��c������F%���x�X���jD�v�2�/�tj~��]����BҶo�*$�_��m�f$���ٗ���y4����H;��hz��R'9�7�pQ����^4��7h��x���< j*Ky��$���3GLWVi��n�����{��^���p��'#ͲL���	diS�4xP�Pu� �Ogf�@��T$���f%y�0��y�/H�]T�Rcd>O;YW;�3�\P�	p�?��UD:�r�>AH���*DOw��o�_ �x{"{\j��6��+�N��C-|��b������[f����v��Nt�:��[���*F}���T�J/���{CP�Q7��1�cO u��bU�S!�=�S.�I������r�T�"�ݽ�t,L�)�Y/nvGKe��Y�����*��E�x �� 5�|gߌ\���k�f�i���M���� �&�a�>���˨I��)��jVYG'�����	>��S�b�d!^����b��v����w�C��ta:�������[^�ikV��Grot���N^Z�(c8c���RQ&�j���"f��r�d��|S����PBE�>������Z��H$��Up�Mb�GиA�(V�pˎ��An:&�Ϗ��R�S譫Ra<���a�g1�� {����q�H���!}Ţ��	��}�K����67:�ؘ�6gm���>��#��|L���R-�OOQR#>��=*H�A�g�����lC��lʸd8�Be#ߐZJR��H"gߊ&�2ń�W A��,�l�7.�_�� �3��;W�^1�WɏIO��jJ6�73~ ��,/����܀�g�S��٩���G�ײ~�g�������c�Yv9�N�;?�uM<%F��������� n��PYYi�q��{�C h��8�kU�h^�����h�s��Zr�pL��=;�b�3'��Y/�'�IR�U)�&M��0�,�ʀW�zD�0c[�I<s�D�>�l�X���� g��TfgG�ϜԒ��d�-.�7c��.D�y�Z��X�|*Ѐ�+�������~���>m$�Xs�H�y�7G3�W��sq7>����0!?�ᐻ�}*�H�T�p��t�M�T�Arq��-0����f���IӓA���;gzj�JxE.�I���?g%y��ЦŨmjB�����1>!D�g�.��`�t TQ
�Z8t7ڽ��T��	o�b���@菳_c��a���~��a�+	B'}�[�KfL��zt��<F�nS��8#�W23��P9�|�]�{��4_�|�З�CJ�1zF����̮@J�ϒٜ\�b�:|
�9g:(g����
�lb�	g�L����І.r�<���i���}P�M,5]^K�>�n[�e�&*�\��o<`��xx�m �(�4��b�b�ә��(�������I*y㉱�Zj��4c�ލJ��`q��y|Sb�k7ռ��5��A�cq�/_�������_�����Y�:�^��sƉ��?��ɾP�P�1�#.�H��uf��� |Va�S}F��A�)�kI55XO��H}�/�К�}F��[�j��qTu%b��Z*8��,���FOQy����LM9�6�{�6�֕��nJ��஻׾�sN�gTX�b/+�s��8`M�̲�l:��:r�����*rm�M=����+��lj�n�;��Å���tY�n�"�۴� ��d��_��\v�9�ȼP���^s���u��±�{J��$�?��q�6�P�2�����$�����*u�;9A���Wӯ���V�[AŦ��j����K�Ɉ�S艥eΜ��LL�$�S܀�������X�㵢��k*�-��[��	4'���V~p�ք���A5S&ֱ�#�h�S�����ͽ�`O{��sd�d�C_��US#����X�UH3VP7��]'�.��~)���Tr7Q��@�"�� �we� (�- G%BLi�h��QWv����Ə�����������hS���\��6�)����B�C��mF�v�8q�[�e�����$�7�7�N9_��6 ���
l޽��H��BZ�mGO��I	VX[~�X�s���e����Cf�H�oò�['����%d��[Wc�Y��.�)��xL67�Ȕ�2�y( ��4���̊0R�R�L�%��\�o�ռ�@��d�J����w5#���<-&�M�c	��ju�����F>��J��S+^����)���R"{�H�s���G���J����������Bx��'�=��x��9Y.��w�B�G�,O�9�*h�� \�o�|M�'��@�_z
�H1��w�k��V���2�8\�J���3fm]gyş��5��W�i�2��F���I���jM���Гʼ��Q�-){v���y(����r=]�7#*l�;�����GL�5��vVBŬ>��CS^��k�:>���(�����d�a�mx��z(�[�cG&V
p4#S�2�D˝s�&�DK�L+CJH	�|-Ȋb�w��D�ݭ�������*'}����v�c����xf7��Yuk ��kM���Ce���ډ,�:�H��1�s���)z��g�r1������GhEl�:d��a�E\�>Y����*��Ǩ��_-=$����A�����,�ְ,'�x�ՃR���`�~�ٌW_f,w�L�#wNޱ\㉀�5bw���d��Nm@D���6W\|l�76{���HsXC�]��Py�?;B"p2�kl�^8����<^�����P�V�)��@��*e�]DA�dR̵g�O\�(8x�����/���),N�v�1�v�O.N��*����k��g��53^ �T9�%ܸ1"'��g����.-����^o�Ԋ��.7?}�����/���z��6��iL)�C��<�"@�my�z�}�TFſC\vgA �8�ha��op�%Y� ��? ��A1�cb����2	�ݽ�MːȌo�΁L��L�*⇓E�A3��~�XȬ홾��
����6�HR#���_�s��Cn&v�d'�� ���w�h�,��所������(_����������w�5n�)S�|7+�n�̇�A�a�`%� ��4.;��Y���[,��	��l�3x�GS ���#nA�Aknة�I��1L)i����@:'�����q:KLU�屨2��w�]��h��G��V�j�VU�OyY��#L�o2,K�h��=ݢ�9���ǅlǅi,�d��
��0o*���ӂj�}>%��L-N���7���gȟ�[�b��0v4��v���x3�kT>w�1q��KǗ)�+$0��7k��m!<Z]���I��S���3m��#�G��ό��l�ܓz{�Emo5����j\o �T[�nO��M��+6����%�5��	�DB�tȼ�N���b$�;DU\9Z�6G�����s"mZ�� ��P~�m�6Q5?cW�T��rq�D�}:qXӞYr�G���=� ��C��k�+����n[H�q�F�P�ǫ	BU36�pB�߅�o�y~�.J�ݠ�C
�V"Ӗ$_A��w�I��$�^��WcXȗ!?��;S+XB0_��kk�M`����B�m�6�!s��߆�x��J�LU��[�f*鲒8�.�Bu��S��^�y���ıaÑ�l��U t���[�4{��[LSd��t�Ǹ���>���H���ڟ�T�='��j K=��:����;2~��U��H�1AQ�U*u5�-ܫ!�G��=�<��������[�E�0�Y)޴�m.�Ů�8�� s�#f�z�ʝ$����uLz(Fdנ0�Q���;a��-����!G ��.�{Z�S}��J���F��5��控�<�q��r�Y\7�5�e�(Ъ�b�64 �Ǫ�]��՝�/2��/48��j��������1���RS�IY�yl��}�!�� ,���������q/��kbGB;���#�ܔv�YO�t%�����o����}�"zJ횜RF�B�QJ��.0]X�:	PQ?6zc21�Եf1�Lѐ�g �����O��%Yp;<U�Dƨ�����~��cH��ߊU<g�T�U���=�i��{�6o��!ފ�㗂��;6E�V^��x�\q0"�<e���¾�$���o�P�m����S���|���kJ���F��cԁ��:��b������钁��{��Uqف���6w���V��<��beb
�T���8�,�R��z�|��I�>��mb�I�����F �h��[ݬ���f8
9��5�����D��3c�|�����'��P,��-���gGX��xٝRΎ	t_�8$s �&%�������c,?K�~F��oYQcp6Q� #�Qq-�M�ua,&���Հ�M��U*_������
f������o�VT���1.z�k��b8��"|6��w �H�2�����M�����\�]��m(���K�M�#綄J��
��^An���K	�%�'��#_� ���T��PjwѺN~o�L��R����[�
�I̲�㈁Te�)��zU��o��욋['�ן7р����z���Y~j��ٔ���T���:%T2vK�L
�"���vz߀v�������J��� OH�r?f�� f0�!�a�H��4w�A�{���{7��
���ti%'���D��S-'�f�B�����0k�t9)b5�x6�zK�2�o<Tل���o^�3��