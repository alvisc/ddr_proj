��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t�������.NT�ɯQ�_�EY�����]|�=�Ăt��@��{D;ӸBr���J��;��?�͠�j\i�ş%m&j��?v�W���tF��NO1���?!T�Tg�U-�(�	Z1��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC. �,"��'��g�	���:)J�U��>F���\(V��S�Y0�$�Sv�ջ'�c�@��mt+�:4�.�Y��X\
��z*WR�||"�i"�����ᓇ!�I+��_�Ph�5�5&ig @���bl����4Lꭱ�jy1Q7�r\X3p �Y|���u	��[e�Ƕ����+Ƴ�K��$[{��ha
����6�{/c�wD��J��R, `�s�K��un�ZOF���_i����T�3��aO�����V���n,R�L���>���
�&c�Qrg!����x�
�%{2�c���'է��7�u��ursf!���͢^�sܻ���@�3���	�����/E�u�T��I�1Q�A��DqH(X1��~^�ۙ�����{���?�k�]d��0��kc���uVB�Q9�?Qw��,�Y�.�zy�6���#�w�q���8��S#q_�E�R ����ɴ6���W$g
ݤШ��d��е_[�1�^OC��o�Ш3U�q��g8�i�#�ugh-M��� ܾ,�T��n���D�w�9���+k��*6���#����ͬ��r\�b@��J�9ϴ���Z�èr���g"d[�\)��0b�M�j�	�ʮP����l���@�����S��g�b�o�[�ki�>Z�O[!ٳ�Ci��j����>�j��</����V��������:�BA%����o���c3�	fe�a�xv♯!F�����FW>��h��鯞Z�=������.��m���>�lE�����٩]F�����A0�0" �F(,Y���$��z���7]#�Q�S��!Z��1��smh��q�&�!�`�T���Z��~�	/�K�$||	�ۖB�?P#���=0[��0="�h83Вr�~���4�?��]�jf�(��cQ�8guŞ�:6�p�TaY<��fYr���a��p��cN���Bz�P!��r@W�`0�19�{�B�2=�?"Kz��Fe����f�^w־��b��HV	MbV,2v�<�i�to�k���7�����5y虢iֹ �ߌ��=If셜���/P�U�Yc��g���~<��k�%�m��u�� �L�i 6�,m�@or@z�ԏ\,��-b~Zk�a7����R�[+�^7�)�	-���;1y>��!��B3�ԓ\��V�!3��b�'rDikC�j`~��/�h&�$^l��,�����RDϔ�f`��==��k�(�3HEJ8�dZ#������ ��^i8��>����+��Tn��C�P���	h q���8�� %^,�&V�4�x�K��50� [�N�1��:��>�L��4-o��9�Z��	���[u �z�r��ۍܬ�Ǥ�=�n�.Ʀ�F����&ޕjśL]���>y�Mа?��Js�6�i�?�~������������7��1��L����*{,�~u͌Z���`\�����f-��'0�:nĴ,�x�d��P��:�R�]����r������H����g�١o�����\J�^��4���MFiy%��.�r[ ��v��!%~�����C�6B��!j��-C'Z=Z�H�Y�yQ�Y[�� �Z�A��R6� �+Q�G�[cqD��p�&r! �O_E ��t��=;o �[�0>@����]GA�$���};��#$vºW�㑢9�I��g<ѳ"X�)�\�$�t�6BU�~�F �%3r��L��$k� �[eLT���y�F����$� ���!Sf�b=��k�5F9��Ս�V�Hi���oyhP���3��U6��8��XJ�[�T,�%U�3*g=�_L9��cE�2��G�J`a��,3�A�Xk�d�ϺHh�(Dd�(BT���X.���-�&Ւ7����to��wp��\g:=z����:����z#�����mܭ$�� �_8����mZ>햃�؜Hf���Z���r�J�[C�WַK.��ʹ��)�-Ū�<!w���f0'@��x��k��-nY� ��>�:�zr�\��� <3BϾ��i{=b�2~y��?	h�C�'8�FU��Й��?���ɐu�8��jk��41'lx��m�e���.�D�'1�(�����-c�yY`3/�����)c�@%�Ў�9'�DF��J%Y�+N[,1����)kD���Q7�[!��� �a��Q�n`2��x���;�@�ix�K*3�=d��:e��j�Ϡdtr^m�,:����:���,zj�� ˣ]�s����v�(�K#�D��@��-SL6`��t�U���t�^t�d,G�>�TИ� <������q���0T�Tܾu<r��ޚ���*��н�#�ˆ^
(#X�G
�����&HtM�Q�Ty#c�J�W�M��W�Zı���"�U A�gDa��$�U�W�-3��r�'�����;�߾7bLXT(��[�Y�E�.�|܍���`�4�oQ3��ݼn g2�^�;���J�.��3ρF$-hl��:����k��M�yB�Ne8C�*(�L����zB�H��9 ����;n��/��h@� �uBG%FH"o�զ�?G���B�0@S{��(%[���h�����ǫܨmϩ��RÌ��!ZT��4]�� �;[�ݾ������0}b��*����W��1b
I�Ԩ}��p������ɉ�r�&q��x��`�O(b,���%p��N]�U�SY^+��5Rˎ�yPep�x�ՂB��ޑ�p��I
eQ�| ��Q\�ֿ�C���[Y|���J���P�g'�.����-H"�u�x�D�/�쬛��ȠE�P'����O�e�����j�S/�d;��ƭe줫��?�%b̛NW��wT9�`�w�5!�Х0�_q�������n�FM�����U��A��__.����ދ�+_�BԾ�Bgd3�Ӕswt��Ћs��~Pi{�Ψ6
S��7Z.� �X?~gf�
�.銫�b�@Bz6�D�_�R�DĤs����څ�>��׎5�W[���S�9��0>-��"h��fŷ���N�Yq�(�)��˨m+���H-@+,N<>i$ം5�_?���N� x}
v�:�N�OC����&Cٌ��P'/�l,��&R;�ư�8���'�%qa��3����	O�M���I��*Z'B�#N�WP!�:f�o��rͪ�.�8�>J�;T�M��9{��@���P�'vy��_	�6���g��)A�y��&���H��K��2�$�_�G��(�q� �S�\��>��EC��ι5q�ř�'�jvMw|dP�z�����^W���ux���~g�\��PY���j6�=aU�SbMX��nn�=m}�a:I�TW�}�A��3�Ā�V=r87�Ύ�
���p%��hz�#^E��\�FZˆe�fC�`{�vp�@H<P���Ź��ž��CH�b��iȄ�mGb�`�8'��Jt��p��a>��N�Ϥ�m�����V�]��u�=G�����ckI'.�e�,�5��8�ruf�� ����QC	حB�����J�g�X��}a�:��6Oj3nZԨ��h��3���v�ٺ��� ���t/?/��><	 g��Xj�jי}QR�`�Je-�4�<���
s��(v��@Jwim�΍��:�&�&��$�MW�������&ݦq���>�����F�P?�M�oK�{B	)�s.$���;�z<����X0p\4b���/k���#
�Uj��e�m��J�
��蛊�xl����|�1L�񗘌;p8|�3��攖���А8
�MSeC̅�v<�q��6�0f󙘙2�D�SSK�35vu�Q��Y���V�,�K�j�Gz���ߢ`:�\�E��k��Iޖ�Ű[o��W�����s=�d(���h�d�&u�U��O!�HzI�d0>�rY^����ԏOܠ�j`� ��9i��ʟε�t'b0oe&��c�}�'�:�{_�yՖ���^P��� O��O﵀��]s{e��ʌ�#(�2�Ӌ�1�,�ܢ�NS��I�1sZ���5f'%�΋P��%C�����8g`K��<j]�U�S~J�Ÿqi�ch�����g�a@;b��b��+H���r�ܔ��{|�5A��ɻvY;�I��u:t0qy&@��k���g�����L�ˡϚ�筯S0&U�̄mp���,KA�$.K�R"VcO�6a$%�+�pc���oA����4o���5A��^�hA�!��|g8`1hs&��L��[�|`Cς��Čiu����<4�i���K8��G�%�bS�=��P�ݘ�vF��O@f����W$�ੁs�h>�zt�->%�i����P��W>Z�S�� ��f9I����Qk�L�7�w���( ų��H��T*�2��W��}�:��^/�?uHV���n��D>ߪ(���/}�2���C�1n�Ȣ̗�3��*6=p��F�'s�<����(��H�QT�(�dZ��^ķ�
�S�M!��6 DqL,�A%�l���]�`�QK��[�R�t�C-@!'ʧ���\ڔ(��p�n��@v�U�<�.���s&�M�r��t+;�i��`CW�uM�1v��Gq�������-䙮Y��Rp^�y��-HK�%c����=ū�26;��r��YS�i��,f��}�%ŗd2�Lז��d]_#x%I�4�˥�`��?7��� 䂂wR��J�X@--�$��B;��O��{��<>�{b�$�++ל≊Z{� �[z�蒚M�r�%df��ew������f����<��@����|�%����9���֮�߼t�0v��k�� ;*��:�+e�8�C�<�U���˼F+C�2i��=:���Yb��ʝ$6�ϒ�K"�U�%w=	aߖ/Xp�LjKo�/ͪ��纫���WiXXl�Ѥ����'���a�
�d;H�ק(� �H=A�aU2�^�2tK��n6>��%�u��-B��b��<�@�)��C�ȟuS8�ǜJl�D�wUk\�|_�At�6&G���18����������4� ��N�4P�םy�t$']��k�SC��\�82����q�..S*N�����T��ᷝ�w���q��VO�E�`�F%��-WR���
�,�6�؉M,QY�A~%u��s�����7�I @>4f�������+a���|���btR�:��dK�-�~���9/;��{�b��!�� ĶW�ןY�"K�)m�1�!��T�@�R�(�у����V��Re/�߻�"�O��|��}Z4��̺��)I�,Oo$��!��De,���(k������[��S��W� �(i���N�����c>{s�F
P<����n�E١�'��͂-}7,�#f�d�e��E��8�*�W�؉s��ԑ8@.��(*�����������q�HR6�8�?x�	*���9@�E�_W�p���"i4��#��]OSY&�����^�2*��p�DƧ���aۏ$\ 7�S��-8��g#.)��a���^j*�.�n累*ǡ:1i������G|���/�]u�4��Sl�"��z�o�$��X ڬAH�AP{�<����=qS���5�*C���X�I��C�d��%V7�v���et�$ �qN�)4�W .�1�����^Ow�WO�'�	Y�x�ؒ,���d=u��ֈQSk�i��Dm~}E�] rhL'�Z̜b*dɂ��kr�����8|��w8��v��{��5�t���(	�o���
:�\?̯�W��F�������]�%;�^�v�g���Pr��%`r�i�׽���JYuZ��t�w���k*���k�ON�t�3ױ}�K�ؚЄ[��@�����tG��tn�@�|6,^�X9��W���_�����\�'f�R��G�?��~��k:��>v��r���B$pA`�_����[�;g�pZuErJb��
��DZ\���7��wxO�\�!�]�V��3��o��=o���#�<�� ij�/7H\�-��)�v�4��B:��h��������k?_�Ǣ٭1󤇟lx��K�����l�����:W���w����K����������m��q-�W�)�E|'FUZ����@��SG��)][�|v��O��(6��eh�[��K�kM]��m!K��<����^������ֆ�ו�0X_#@t99ql3����>����E�X7~		�Y�����1�V1H,6P����5dg8��O�	����([����g��$Q=���
�Xb}�o�(Y
{��3����ݟf�g<����8�nk�7���a�h1�f����p�jy{�	�W6�Y�?�p�DB�剩C��a����(D�k�\��{�0���y8�����XF�r֕FKၻ���<���}�$�	ag��n�N��m��$�r��LF��C����Ks��j��68c��7�z�Ի�Դ,�	�������D̛��T��r�n堧����8,{��M����}٫!SfmaS���cJlA��]�+��ߪ���\� ���R0_s�ՠ�7�pQkn���zV�_�^�ρ�> �o+jh�CSξ2A4bG>v�$��t�d�%��v2��Ď�t[� $�ח�:��9qP�m�@j�*��i����~ys� �p�w,+��Y��h���֚ҽ��p�=�T�Q����r�m�'9��Rژę�߈vEE�V�.wa�.�.0{��qV�%��]��m�stH�v-p��)-�:����U���μl�uS��X���/�o�ٹ�G�,�<�T�����-�v�/!ƫ�$��%5����D��.�`䆲�M&��D#QG��=%/i��R4i�O7�͟�Ӽ�K�G:q��l4/b��x�A�)�����r�(0lx�d5�c#~�T���ʲ�P��c��Kl�����Q
/(���� ,�E=Q�9�vǖZ��u��,_���b�U#��t�J�V��h�z=Q7*�����P��� k�!�^��w�iq
^����z�q�����䓳�o���t�y�.�0���J4\��V%�D3�H:	U�"_�����?�����@��y\	7$xN*?��8���p435�^�wJ�2���uv��cq�X�eUY9��K��#/��#���_,O��na�������(�X�!Xj���m�90:�X�N���
�h��`�ِ��cx��֒��YsY#�i��>܀ķb�VJ ���˃�n����4{���a�|�M���oи'NgNXyYvH�Z�E�vW '��R�pW[�@��B���� f�w���}�V�$�sʧ��%͍#4�pG��S�E�� ����`Yұ'3��n����/���k�OQ�g���V����2+��)R����#��mn��R�{]a�\'BH��z;�_�p���E֪1�`�H1@7s��%�:��
�dR�MJ����[�,X��X�0��m�G6M�H�t��9b6�B�&n�?�HT��p���R ��z�;P��&OE��e=�c'�J�lG$�aC��qپ������K7�*M�21Lj��YW��D�_ �⁀�.5F�=u@́�ݽrW�*`U�=��R28=���+K��O�RRZh$L3A�1=?�BA,yC35�yv	8pO�z2_w��Y��z�9������z�����m����u�.�#�3�fI{�SZ)eJZ���a��|z�7��4���-�U5�1����m�c�Kx0���116|�(�����"��QWd�����Ή/�L��#d��'֐P/?=��#Փg^r#\<ͅeq�����k�-��
���TN�$Q[�QJ~X��ԇ�*��U��{��墦u2/��A�7x&�B����/���#pH�;l#��S`7��І�zt����SNӈ>J:�O3�|�UQ���Q����/Rk���xl��y�m��rZ+:�	���n�H�"8�e�`6o�w���j��<�V}�ho��a� �^5c0ޕ�[�Qw��vU4.��EҲ'�}H6�����n���=�b}:D�������^���ӴKLv��jn��ao�	��)q�ܸz`ymz�^؛}ԬՆ�7YdX�%jd������!D���v�T��y���06�;����Ԫ��O-t�6��V$z���>A��;��O\�;�e�au�)�1,0��V�@����:�9������򯵢8nZC����~�O������C�L��*oVw2��?a�xI�� 4o@rmZK=����3�\2��2��'P�H`�k'�WI*���궷�n��	jZ����VLc�={ڡ�0P���ؔ�^繻���OƎu_*���+�Hуa�wd��vTWr
�X�	B��S�I;�XZ{���:�t`���P�phV�T�F��Q�u�:O�C����*wv�b*4���V>V�N�|��N�J�an����h�|C[�F�
�<A"�TMm�E�X�G��0��<�Ӑ&�g6u�|Uӳ�\�o�3�uf���ZhU<#��mZi��� 
�T�5�}�Og!cNI̷$����S�v�S�wb[���1�C���B�)(���'����߆]1MG��{Y�n��7O/�e�6-X3�VJ�x'��˼7��>���c�gB�+^��%m��H��n���P�-��M�x&�<��V$ƲW$�jD����J�}���'�����;�ih(vɛɫ\�D��i�d&�xꊚC�W�j�����j�qCC�̹�b�'*��SI��Êv)���$�y$���)^l�Q,�|���1��CR�ҝn{��J����XR�hf2��/�: _�[C�,�&��H�?�������fs�?����S��O���E_e�2P���Q�q����GGi�o������<�LZ�*���x�bS��0��	m�ֈ�)[�����L�X�Q�G����qa$ܤ�[���6e����� ��_ʗ_x̄��������O`��H��Kg����pYܮd�qt{'H�D����6#� �r�`�h9q�f!8��9V�:4�Ǖ}yW���ʥ�T��,1����Id5*��i�����91<��9�+�f�ay.��L%�,�훴���N�b���P�&�Ia�&�R�Sj ��F��ψ)�1$�Q��Z�i9HI���\_p����O��e�4�	|7c	�0�z;�v�x
�~�§���W��hbu[�#����;Z۰(:��@���#\^�A@3wܝ:B�ۯ�� �<.4C�#r����ua��Ge�N��I.r9�JaR-:�vp�Yr9�<��y���El�RgoR��Fd��^���9���(���8��[L���3�g�	P���l��w�J��wuӛ(�b���x��+!��)�M�_�Ԥ s�����Y���3�\~_3Q�J��Ekr�6�4�C��>
yQ�����G��o��8hgv�0���).4� Q��]���P��n��.���-��,��X*��:x�놜�*i�-�h��7��Kl��{b��T�=� ��g�@>R��g(�$�g�ⶁq�Y�Ǐ���ĞY���?�"ߍ��%>-[��
�O����ح�{ļG�K�'\�U��� �e�9{c9�,�G��4S+��'<z�wd��]�c�_��օ�-�pZa[!u���pԩ��v*I�˭Y�6ԛb:e�-��W&��Ǉ�P� ��i�8N����K�ˉ�q��nI�UN�aG�q�rn���@c���A�ʬ3��s�;c;e2mcCw;��열~!��$�^�-ic����TN9(3g��Z']��%��D���,cW�[�!LVZ��}�N*�� �ڂVLoiPUB�q���9h���ӫZQ�����P�֙��C[|���ġZ�?��x���5�P���~���6kW�R��ͮ�g�b��V�d��E�@�q�m���I�V�CI/���'�f,Xw�Ð�� ��a ��XY7�D`;$���$�a)�T��I��a�f��X�q�1E���LVӟ��i۞��`_'��A����4I6�3��ta
�B�ɔi-x^�c9��Db�)�B�-ˇ��A
�eI� MY�&��t���d!��HH���&�#k}�޽d��٢�Ƨ�� =xR�Kٰ������*Ή�d��y�۟~�x�0[��-�|"P(�j����S�9T&�\����3��W�_��W�NY�G��Ń�I%(2�r�+�p�L�s:��2z(p� l}��1��k�Im�71���SR0�O}�ߍnY����>����S�3։��#���䋓�o�.)b����ŊC���uGX������q��A�"���+��}J0��ǰ���k���J/S�y��+����;y������ }SDB1���{�sj0�ZG���JfGv�|�O~2��O4Q	y����z���N�i�z��-H���V����eu�K�ڒ�C0�G�u~,�30[�1^ց�j�-�+�lGib:~����sA ��e"L�\��Wi�ogHW�V�����P��y���"�g%��<�2r|�IN^��"[a�(��}F���&y�{�,ͥa�AS�.>;TE�j��T~q^~�Ow�dT1�ף��`��E���Ë�i$�?&B�?�AkdE�{/k����3B*�4�T�܆����YBCԼl��|�጗M/�[�D����K?+�)���hcS1�)��TN�{�R�n����h_�(C���c�A\�9Hۖ>�`Ϫ_uR�߿�\�`�R����0ٜ�9�4{�����|%��'�t���\��Y�Gi�h���!��F0Q�mU4n]_bl�V�C�nh�Ղ��3�c�ތG2�!Y��\-19�]�����,k�Xs$��Y�f�o?@&�Y���M��Z�h̓Ɨ�7�J����ޔ�`��W���q�$���8�M�5�C�v�R}�����G��rxp�3��!6k�s|C��W�!�-	�O�jT%d�>�/\���1��\#2PnH�d�����`�Q��-�M}�[�S�9��c����A�#��]TL��@�%ɍ��9-��ģ���2a#����Z�N/LB3�^ �Uz{�PZX����jv������Qby�K�B����NB �^�c���mOl�s�:��8�c+�:���4}�<<��]"5T�Ϊ���w>)m !�G'*K�b ,��i���9�0�xR��dwu<l%ڵ� c����*�����eA�bddw��k���Q���^
���<�i���8��'�f�q��{27��-�j#�.�2!��TL��(��;F�;*KJr��*�z�Z�7��־A0� �ӐV�ݨ=gmO�r,d��j���fI�e�:��p��'.Ex|�� )0�9���nT����Ey�V2�������|�RrxzL��?l