��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t�������.NT�ɯQ�_�EY�����]|�=�Ăt��@��{D;ӸBr���J��;��?�͠�j\i�ş%m&j��?v�W���tF��NO1���?!T�Tg�U-�(�	Z1��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC. �,"��'��g�	���:)J�U��>F���\(V��S�Y0�$�Sv�ջ'�c�@��mt+�:4�.�Y��X\
��z*WR�||"�i"�����ᓇ!�I+��_�Ph�5�5&ig @���bl����4Lꭱ�jy1Q7�r\X3p �Y|���u	��[e�Ƕ����+Ƴ�K��$[{��ha
����6�{/c�wD��J��R, `�s�K+Ke%G���N�;5LR��>7���F�dR�;�#a�=�?�c�=m#����?�5�^���f+ns�����
��%p�2�P��}��'!*b�6�H��V%wX��oܲ���|9�F >��T��ކ)f�`q��'����O:��u�-����Z:�eN�[��d����.}[�S�H����o8Z�e�� a�]���W�JU����m�G�E�L���4�$�V����x��(V�&N�%.򔨖.q��$���ĈOKP��*�`�ź����v�c�^���i��FGI��Sr�x���p&w���.�s�Q_z�'�.Ӎ�u�j^y�5�&����H�v9���MX��Ms]!o�]8�/>@SE�X�fxf��R�T�@F�׽ϊ'O�U�[��^�������b�q��<��T�a���`�0���
U��g�ZY���	�1�g�vI�M�����L�#���i�ч���J#֌�#j��g!�_*�[D�	��4�ǆ��#A�<�֚�q�Q��;�a�??/��6�1�5���]��V���Y4N!~���A�6mFM2�Ҧ?^�Q6��}����R�Z�^�!��YdW(�uRN�P�R�Q���i��(����֞��.�p�,ƠaS�La�ԯ�q���A���Zp�?v ,)�jb3Y�8|A��v�����8z�q�VK�_��z��6��f�W��d���6������m����~>�W!�8'l�/bU�z
�Hq|��0K!��3VT�{Uv	��{��2w~�z�̫p.�:���K� ��х�a=U���q���x��]�1�,�HKr�F���x��P�����?��&L�JNB˹�Q�r�Jj�l{<-�!qʕD���U@Z��G�B����>X�7�.�sh:�r�	��J �m)�����!��Ǳ��bNܱ�E�EW}�R� �&��؆���܊��:�P���)�6�����E'��7��[�O�'5b"/X����,��d�*v��d�c�������E�8����n�p�j���y��+�H"����i�s�.M��
։��/�@ob0�;k#�^24�2'q[������8���|�K�0G�QődCƶ�TG>�T�̷$A}UT_ٸ�(H��z�V̊�0��S�2�+-PGAZl�sb���������
"��:���h�	=���*dp�;��^�9��G*.6'E�����l���\��  $}�{��sϘ�Z����:�*���Ea�),X�n�ٷ��FX7ռ��o��$�	~>��킂S�qRս�Y�L�@f�Jy��� �����Ў�ڷ���Ù���ʗn8Ow�G�&��I��8�X�υG]���E�mYu*��F��O�N�.ie��ه78G�(}�rY�@�t� �6`���2g���Zep���a3�q��{��帝�X��7*�\b��S��x�߄ɳ���WV�7�LI���G�S��~��8 [C��L���5U�h�-��2�i�>�ˎSc��Wg��.
�ؾ}���.M�((\B�r��ਜ��������8rBX���,c�}�]�*�q@~ZI�M͒�P�i�M���?�
�0۬�H�^M>�f�UIJB�`'�jm2B腭c
8�+�*kj4bjut]�ls ٽ����n:����^�Pq��xli)!+�{�	�2�[nmQaN�-Y�:�S�`��.�"�)�{������y���-���Z���;��IB�3���zO,?�Y�����h��{��S�@NJ^���~��q��������]J��z`�f��d]��ó�G�p?ʝG&����c\(e�nVʑei��3��7r�h��>�WiqKr@A�S�wEV\�Չ������L�7�������f�豧Ù���}�˶Nr|يg��'��{WWo�z�e Q�y��'�k��.��';��l���Š{�VX, +y(�]����i�q�\�QX�~�.�2Ũ�l��� E2�?[R�v��0�o�����]�{�ԑG�sǼr���"\Ҿi�[�
@��oTw����mY{̯ę� ;8��,�Z���Ì�D��̶:�u��i%��c�`M	W���Ak���@s��}A>So��M��ڂJ��mak+j���j}x{��wz ����\t��̬d88��j�HQ�_2�02��y���#���-e�8k�@����H�T�o;Ⱥ�}��Id����p�}*��ݻ~�%L7�8">�����l�^�?�Zc^��U]IM\�~\;���Z�����m�uq�=3�^�,��ӏ��	��\a}�2W���2���z¿pu]�Z��rE��So��CZ2=��bj��_fE�$Ku ����w�j���^��̾.t����5�_o�����#����v`E��7�j����Z��HG���)��-��|.����2j���bF�r��!�b��.o���k�}�6�Ճ���l�K$��4�,ѹ�{���J���nT���"�b�U�d�_N�7��a�܈�ʵ�c�0���?R+�UBT�s����E�>�&l�Ĉ���-�ޤF��J���Hf7`D�z�h7��a6�[*IW٠3��<D`�Cը�]{(ϫY%��$�r��{��67U��8�g$q��jU4�[���Z$\�����+���{�S���L7���ϵg���
��B�~:&6`�_�㤚�a�`:/4���r���h�_#K�Ҙ��{}`k};��g[BP�}�Ů
ަ�]4��п}�\=����i�:��ޡ��B(��2WM0e�g5Q���Re���D n}�L"�Ǌs�
����D^?��n�WS׎���<V@�kn%s %�؂}���Ύ	��qG�n[SM���p��}u3�R�:n��qx���g	�E�Y�G��	e���'��_�e�x��a�~�?���f^b$׌��:�tp��]�����v:rf� 1�g8)U͍�2�I���P/b��|��QJ��z�h��z���Ր$���3�߂�(�r7���{y��&7���?>���wx��V����ޒ}�o��ވ
�,C����:�
6�{|z=��l��SC횒C���S��3���]�� *�p�i8F��U�[�R����:48�E5�l r
`UjV3ێ��:�twno�,*ߕ#��n��"&욮��~&�__}HG����鮢��I�X��#�}���!�TA�9m�|��y��$x��|�q��Eax�cIs�J�G�.׹����v=�hY�]r�� E'"��$x��Ď�4���NXˉ�kLe��:,�LܑT]5v{8R$�A��>|'�����~���ͼ��X�3�o�}�i'��]���}�(ZqN@kIa}�
1w˯U�-e�^~���e�:�8�֏^��ͪmQX��� �X�����~�^5�Wj,pų�����,ML�d8~�]�iY�3�`5��_۹86�j�N
�J�r�wFHH�m��Hb%d�=��Q]h�ت	iO0�� �==��>U��RbPZ��yԐ���5@w�������Mc%�s��5�c�?0�m������G��DmdZ��3���g�*�+�P;��k�c���P;�=�6Ŵ� tu:�K�f�������i�U���E�V15n(��
E�hOy����@�-�����T
r>������U5����:Yܦ��`�Y�;i��w�6N�!���eh������KZ�dJ�e��M*�󙠬z�h�E/�<�)��l����lD�t8�d�(������xu.'y��zA�I8
=�W??p3
%�?^�Bޯ1�Д+Bټ�uf�aCC 8�@�<¸��]E���]2x����C�4���=�l�C�Ʃ����"�XS+~\�U'�]���J��V�q�P�vmZ�w=&O����( s�X1�K����Y6=h�j�@�!xU���l_
G_;�=7��Q�h ��`@�p!ZD��
�0#�9��D?��99�[���?�R�~@ 7��ἓ�&�#Ld�! ����yCG<N%���C	�dD�|�Q7z����E����ҧ�SW@\�6z A��v�P0�җ������ċt�'�xF�?Κ�'�j�EG0i�n��X��ԭ=2E��RE�pA�	��&��*G�O+�dg��B���#�4�ک�>���V*o��r�}�և�4o���9:�5L��.�<�Mwξ�ޤt0.�m�ٙ�q
SU�E�\�
_��RaEO;�U��|J��~�F�Mj͹*K�Q�q �Z�aH8��`�3l�w&�z6�������e��0�[.Ni�/)"�_"'�TM�Hiq�/N�_��#\�S��q�/s|D��53�>M�ҼL�H�0(%�5���ڱ��8ӈ���rD���#a;w1
>a��)
�n�?�2���&ޕ_!�Gb��K��w�+n �-%3REu�td�1�詰�!��I�s�L���B����K�F�;��;�T~^)�<�əh8ݍ�|!�1fi5�*�b�����:7�ktp���JfDe���5f��|F��+ΌYgX$4"a@�:��g�i{C�IR���G������[%!�X?U�_�_yņ2�V�F����M�A���`J��(�ב ���g%<r��T��ֽn&Z|-�w�*֏t��:�?6evȋ�"u�=�� ��mB)<�u؇����m.���?��8XB����k��8,E*e��|Ƨ�$W߿˛��vI���X�0������q�}���!-��t��I��L���4ڇ�4�����ׄ�K�މ=�@�I� v�^!('�oh��*)iyl�,�|�l���}�(�%��J��5
B<9�"G�"��	��AS���a�@�(���� ����7���j:�5f��0�|P�ؕgc-2��a������S��2����J�Qc�K�q:d-{�\�Ë�sH�9�f��>��L�o�
��֮A��[����å[�g�!��XS�ȓh̖���I:��cFB�t�Z.<?