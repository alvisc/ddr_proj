��/  ?)��ݟJ�9�����Nm��X�[�`�������A-A}�٨�p�[̼_;R��RX��8FV�5�����E��m�O���ő���p:��iT��� 	$Py�#�l�r4rVs��l%0"8����hZe���EΒ!��#��Ɇ�>�h<�����:<�)��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HCZ�C�Ru�����[H��22P^��{������6�a�WN8�L�u�E�>F5��o{�R~�Y\m�Ȕ.��K�Q�ց2.����/8��cG��B�+�%Y栠��'ޭ�--j��7��ml.���~j�n����©�kh�ؐ��=?�^J.W�Ս�8�"n�B,�U��,�qQ�0��'vI�?�֐`6^�fv����x�Bڻ�.8��9X\�7������TиEm�;����ME`���͎�ݱ�tĳ�U�����Qw�_� �6Тj�&[+�{˲
���Vŋ3`��9b�ϡ<|�9 L�p����\�%p�+aNߎ��l�;�0�)��Q�؍a5O<�8k�P��gM5�5�+}���?�h��ᤊ7d?4��_ڼ������E)�N˴vUK���Z1����)�?�APB�7���p����-DҨ���DV+Vy��3��R��T��E���sǊ�����j���JD#���!����C�Ʋ#�+H�6�8s��s]kFO_҈��r�b�L�* X�+Ƚ�b�V�P��E�2A��%�5n�	���l�#4\��B����?"ʕ����4@e�y��loa4#��z�hM��y(��3�贶�)�Mű� ��$G���I�f
)U�Khg�-4	)&I;�Ť�c ��!��n���?w�q�O#Y1�b9�x�bub�I�4Z��?E*T��9������#�W����#'��_�T=0>-G�{��j��U�O��8��5���J��t�/����=I��|��D3�T�4�$;8,��Ç�#Qk.QwdC���ш���MV�":��3�$���Q�,�=�ѹ4����U�n�A����K�6�#V�����|�kq镐�ӿjI#����@�^tgm��]�42D�+|}�
�G	�q�eR���G���I"08Ƹ�!J���8:C0���޽�i��_��cWB�� �����\O��㣔Rw_��"�ƳMX�8�Ҭʤ�5q�f͔/5u��\��7%�t>��������߆`m���P<�@�r����� �[�j���u�ܚ1��,�ѻ��d.RZ�m)��JMEQ�3*������EV���Ǜ�*1����|��&�3UY��5�e���_[]��h�ن��)�M6=����+�r�^����CE�%��>pu}S�g�g�������eo*�+�"%�����L�m-?�R����K���W�&�2d4x�����\����7C���`?O���L~�����ш.�#l�[+>�;I����s�9�+n��C�́�O�vc�� jC��!�6�"��,�gP��8�R�����5����`�{���M*��Po�I;03P��"��^�#mr��moF$a�9�!��
�ۂIP�#;�Y7)"X�c�3���c�.B�e�=^���`�1�W��#fЮL��N�fڟ�";�����P����B�Vb�ʑ�ni��c�X����f�8Ș���Z�[�4N�)�υ�<R���wʷ���R[Ϳ���(�^��lc�����6!]�{*��e�T�}O�ʎ��i,s��υذ~���!�:�<6�m���&B�ف�s��Ł"�>�\�n9+ؾ%0��t�}��fsJ��T�|���~l0_�[
k�_��ַ�,�ĿTא���/A�/��A��L^��=zs莰@i
�o�&�W�X�G҆�{Ԩ����ȩ=�WO�&�m�̈́�m+�e�a����'� X-~��/A/13�:�ʩ2�L�N����sA���|(p�}���%��WS!\�������� !���d�6���(�H�h��Y�Vj��Y�:_����n$�>����j˺	c�V�&a۪���Ap�A%�r 6�Q�����L����hX��������wS�'�ع���}l��.Ȗ��*���CI)����g�r�kSۥ�Y�E^��L���uZS���Վ}�%�����150��!'9�	�T���P�=)=,4��R&��{��JPp��u��9D�"�&8��Cr;mX�X^�_�>ͬc#?p Y��:g�S�� Q� �~�N&��֍+�`�X�Ӕ�
6�+�W�_7h*�ň� ��Ҧc��|�jv	������+���D�*�6v3��ɚm2;��;�$�;C*Rg��@E�Y�c�$��&йlA����I�G����f
Q҅w�O��!�w��	�n{�>gjS�jx��P������F�b�擩��
��o$�����d3exVb����+�޺���� loZDܵd4�7oMaa�Zk��<�p/�wC��<��
����;�+Hl܀t���W���N�5�_�
{�җ���p�u���_IS�C��G�ߗU��^HYu��u�O��̿��6�t�1��@k�A#{W_�]ʌ%d-�R�2^'ȍ��{G��5�ÙT���9�
��G�)���-L[�qr�������5uy�'H\&P��t���4s�,�ǎ����Q����K ^5�9��,"%���^Z]rGn����,�ʄy{�C��&:�/�#�û��^" ��6u��6K�^�C��t��9�"��}����{�}��,J��a=F<��
�0�8scɲ�  ͇S�O��?��"?|?�
+<�C��Dzk�K��m��1�+��b	�T�+��}f<A�Oi�C�e����f��`�ꖑ�8�۲��S��ⱆ��r�^&xѾ��E��	��]���Fo_z:k��$�Ed�.|�f���3�^�����딱}+� ��jm��jۤ�WN�V	���K�^F��tC���3����ֱv��\	b~h��]�N���������o����E[�c��3Wu�on�3\("�����ў�r�nP����YE>T �g��<Z���];8�!+�[)W&?2�cyI�]{��1��Y�������0�����+�T"	��&���Gɛ4B<�z�@V�#�W���=|�6��4�c��[��U���&�9���YHH8�!���Ɯ�0?f^�F�v/�?#aP�vGbʭ=�_o�Uv��1",��i�z֑�>�4R�i^,��8������`F_�ΰ2���r�(D�ujn�Zͷ�/�J	J��^7)���3i�:uU����@e �=Ld}��B�N��'ŃC_Sr�S�J�H�X.s/T�,~a�H+��ֆ�W.X��o��*�S�� ��ؙnW���ے;/X�0��Ù�RI��Jy+I�__"M�\E=�p��e��?ƺ�6Y�ݰ���A�� �OPI�r2�nh�����{޵�y@Уr�-òtL��~orJ�ײ'`��E`��NB,X�bg�
����,���$���=����Ue�������H���Y���1@"��/��ˆکw�*`��EL�[5�g�^3��V$]���۳N��Pͅ�Sڶ��/<�� hn�`����b�3���S�G��'�"�z�S�kư�w��¹J�C����g��.!湉K8N�����*����p�=;�({���E�L��sRM�~�Ƭ��2��k ��6I�7��ˣW�5��^�GWi��/���w��!�<!In���T��_�Am�u�^l���]���];0aAㆰ�����a���	�1e[7x��gVz��W��
�1��W�J�Q1�)�G
�
��9�����]`�������0F�T��y��� �<U����5���Z���?q�v>�Xۣ >��Dt��Y�J��6�϶wt���p��t��^��[���[���Y������N��D��#�[�ŷ� �UL��\�%����W3����`f�=�w��P�b2�-ʹ;��V�BTJG,��� �d�J/�=d�Q@2�� B���B������cb�s��o�R�d��{No:o�o��U��Җ~q;,�'��Tȧ��m[��w�k<�f�^��{Z��]C�Gg5�)�v�0b;qh�aa� �0?)sse��'�gq�0s?3�z�C;�nnW����G�/�o�!>���k`Ws�e��,��x�M��Z�}��R/���/�_j8,����l����>U��k;�qʐ����6T!� ��}��]���V�Nf/�,��d���%P_I��V�SN�_3�\�1ٿ�q��A2�ђZ��8U��{L�ce�@�Ž&��y�*#F���Wr@󛜰{����/�A^�6��~��}�b�����?�ML�c�[�NB�2B��a��a\*�T���k�T�wt+��tsm�l<�Z,ҠLO��?�$�0��¬ZځiC�rYg:	@ ��	��X?@�Dj� ׈W�z|U�EP����?؄�Q��H��A��E��t���1mO���2s��-���54v;���[���	C� 2=Ŗ�\`��wK�=��D�U.1�Oa���f��c��0RXn��˙"I[0mzc�ɏ�0Y\)��F�zT)1�nѬ��d��0P�3���t��Gค����
B�ÛI�2|{�|VA�X�OV;��+y{`)��Dp__Vt8K�ok.�4�&9����D����x�f�/�D��K��DrŽM��1�~f��ë[��-�oY�Z���js�J�S&�s�����L�0�H�[��ڝ~u� ��h��ݺ�+��/{�W�P�,<��nC��K	����]۶��sè��`%��i3�F�h��
Ǣf`e�F�	�7�H�a!�-�����{BS�S���9�D��P�6�k�Ȯ0�-�k��鮼�b�f�1߰D~#Q �A�l��`+vjgV�C<�J���؛�p>��`���@�����=�ٛ
���2ğ�D��Q_�����%<^����siY�RV��Վ�?x�/�_��
���\)��4��}u*��c�:��M�*�ɜ3����x#��͗��~N�Sb�iz�H|*�4�&=ۈ���Y���Q��l�iEA|���
�D��U��BU"�}��W0���:�'�5��tA�	�^���A�k$���L[����JÅQ��u=�c��w�39C��VUG52o�"�e��&�1�D�L%��^kH�X�e�;3!����;~��]'����:GȠ#��:瞠+���[��'�l����G��!�a�D[P�񶯯� k^ָ;>L�	�T��W�;�2�LMj�A��5Pq��V����G��Ww���k�Y
t����+yF�ly`���/��=�j�7țR{�a���B��+5�����1l�$���+%��`X�G���M��a#O��V��C�<�퐬yrD���m-�H���5�����4��|�h��pWk/��&\%�FF�F�3���G(�\��
qP��7$i�E�5>�ĳ��C;�����[Ѱ�9#���{
sA��F����j��o��fa�4���R��2�Eb��y�M6#8�-���0�`���p�Öx�1B?���_�Yٸ��TD����{R;��w[-\�p�p�\�'%I�NK3{8��"�L�L�3$1E꾧n�§Oǅd��s�۰Z6��XQ������'E�<c�2�{���f:FP1�E?q�9)H�5w�gc3!���鮱��P�g����A�Y���6%O̡~����|�(0�w ;-����%b֛I���zgH�M��U��E<5�&p�0���Wt��K;q��~�o7F��w0�c9�<��^�)����Ҕ��Dj��&�<����w[��37�k/ƒ9�z3'C>�{{,~�J/��2��[a����|�i� ��M^�U�)ݧf�m7`ϮOeǝRw�mN�f1����Ïj�	ڽ�M2ǹWe�_��d h��:CI����}M��C����B/Mr֡���r���eV�h�?��h�oC���y���O����Db27h�wa���`�~�.q��A� jyD*�\�W�߱��}l�,�y�>!�w�:[��=fփV�bU[����&�t�e�$!]׻���B�MxzsOеxk�C�G~K?����R�V�E�ҍh#�1c��� W�h�e˄�l��|�X�nbf �F�|��y	���ݍeL��\oU���`�+F;n���/����ԯ��?��B]�SU�y�-�tE���?)qgN(m�Nnڐ\RL�n�۫ݯ���IjP`�����s�ރ���5 �����vW��t�z�ԑ}ÖCy=f�&�����K';xQ1�/���̮�۸�h�(��fj_`=V��V{�N�&J�%`:v2�:��G
9��.ԋ�	^Rް�@)_��[M���x,�(�������t������>B�k@+�ڼfefF3|e���I�z_+�W�^�����g˟���>wB�D� ?eC3�ǀ�^U��a��U�9�9�n��c�)�C��B��W뱳��Q�Q�Xapi�`|���B*����m `�����*�D���&SU�	�'�O�B�$hP|�k��ӖHd��R�֋֦��C�IK1�V,��_�>�m揵{/Y�މc��JDe�a5��µ���D~�*���XZ&��5Â�U[�`�-�(���"�Q�%S��6���~�eqO�U���s l�Vń��K��T��]�?�${PTP���Q��{j�n==�@�^wP��+j|G���!{{W����jWQih�g��m�>JЯL�o7���)5Q�C%r�&����?�,x}H_Q�R?�	ý��	���2�C��{O���Q�t����35ܯ�w��9ũ���:�#I�6��'�i��`U��X�iK(q���sC��W�Q�t	E��`���Ib�lJ`��^|���0B:���ި2-2�W�c��V^(���bH���n����1�/����I>]e��.+=����u�@�gX��&(
����NSx���f��q�ޙB�b�W���:e#�3(�Z���𠒦��2L~	,�,�q�m��k�5�0�o��4���`9���`Co��[�~��E����b|ʯo~U�)�*�	����p�e�oA�㷄��e���/JL는�[��վ���������`���_�g���n�[��#ò��p��^���GamI�oRp��\����X��.��I�_S���^c����w���u2ͽ���N#5�Ꙅq�r����ˍY+�D���ױ��m�*����A/�$f�<���
�Im\rF�q�=�p�Y��r��`͑��Ǽݹ��U&���R��ҏA&���݀[�\D��"�`�k�e��N�����|��3���4�  ���"�a�i��'��{i$�1����K3�D���k�ǩnYt)e��my��{�����ʌ��Ǩ���5Y���"u8_�4�wv��Xlc_�����)��o�k��-�]�զ�4�6;�4���I�1��!�u �r��M���c�/����_sWs��DEG��ꏰ��o��^/$`nc�r.5��	���^����񧒈r}.M�������f^g����\vu5�|�Ss������K��.'� �'jG�@Ƞ?��R���'� �/�T<{�Z��vt5�͚ZA7q������@�L��{W���^(C�jS�#��VG$�ͨn�<�{������:$�-l?�5	�� ͧi���h�Q�I��/Jt ���e���(]�F��Sw}t���(37��}����t�Y)����u��R�H�[�"���˥[�o���I�ǩ������x!2N5p���S�ZU3vݦ�vgh�G��3��d���v%���Q�)�w��'9�Vx)�V���;�δ�_j'ظ�#Uؿ"8+UsUۆ�	� �P΁{]��-�Je�76<\k��ڷ�i��쬕"�V�BZ{�$�42P|����'��]L�@�A�5϶��Gف^�)�"ܦ!��]E�
�G�`��˘�mੱU��p������@Uw�%Ѡ�ņ��hﵕ��h��d�m�C���Կ�T�9�����=�(�X�R�f��,��/���!ꓧr]@��[�N��׀Mt3~I�����+ 5Og�����O���0m J� ���Q��k�QK�&^�����^rk�s���C��`=0]0O?C,�!�ۍ� r�1��
�d��'x%J�AFI�/�X�F^���@z9c��D�T��BZ�w����kb��$�� ��Mט�/�Iy�E��@����&���L�H,C�y!l60�-ݪy��_���z-@���Z��t �,h�:��x	��SB޺�.�6Q���b_�i���iս���Ol���a7&�6��]�x�
v���dX��į�
Ta*K6(�W��%3�a]��?(õ�vp����\B4f7�d�/e%��U�<f?)��:�{�m���D��N�'8����Y����r�A%�S��H���;j��q��C���"����}Dٟ��h�@j��A�6%S���R����%$� �u	ہL�-F�5��L"�z�
*6�2V]F�+/�TP��g�W��[-�����xs?g���F�AM�G��u�����q��&�|��K�,<�~DH�Y�4-����J�����>��Ō��= ����$��4����p2�O6�[
��w}����j�P���E��I�YZ�\��@w�� r,���Jy1ʀwJ�ѥ�s��L=ZR4��jna1y�	z��Oꍀ�2��+Z����̔՚Z� ��|O�"��b1[юTIQs��q�s�me{?�'t!`{ej�Rj*G��2X�(A5�]�E
��~��|a���Qlzew���lϩ��9��ђQ�H��Fd�{صq�yDJ}�����.[�t�R48�XM���}=�1�uga�L����/��Y81e*�˂ԝ��d���)E,��vB�V��tW�h��O��W��8��2��͗Ƌ;�d��2C5�Mz�l�w����̾��U'+�cF�l�o�5Y���LG�N:m�47��N�*����Ƈl��r
�fhL;V���ެ��<�^�>>��2F��7�6D��L!qa�+/ުW�x�F����f�Zc��D3���E=6�R�8�>pc�_��;��2���,Dk��G$�f��E}zJ˷g=�E�J�-���tP�.�c�^��%�:�vwZ�>gB�����B�>w��a�&�u�������1Ґ�]z��|4sz�#_ж
ֱ��R���>ۋ@P~�e����lZ�m���h �F��o�	��~�Y��R�����C����s+^u�N.�/�U��|��K��%U������=/Lnm"�p�dA�R 5#�}��8dTY��u]u ��E>~cv��1���?�dlnKu_*{�t�f��V�D�u�B�/���	��v�Ax���O��v�v�����"8ԍ�Qc�<�Q�ڦ)=����fI6��GaԂ>:C�ݡ�pW�~jx��R1V�T(�u��h��_���� >�]���{ҽ�% d�D�p���Xܱ�u������Yz���������������G�$�m��O���j����~�?c':v�0I��Ȃ�VHLBۿ�j�2�����H⣌kY|F �ĕ�M��90�§��"7�3��Z+9���N�g�#��Yw�?U��$C{��P��3�i��(�(\?�?�M���`�U>|�����%e���Qv����V"������fpkv��'��#�\��Tz��Ӗx+���Q���o���K�뼵a�B%|�x����M���Os�
��HV'��&|*y�b����;�A���w:�ܗ��s^�/_���q��[?X����Ә�Ǟ7�۴7&yZg(찻A7����"E
(N�-eQ�}�0��H0vvR���#]�$��sP%�΀��/��������z�:Ml�	A�}���a���;�����TQ�:�����7��� �6a��@����l_��<�M�C�9t ��h{LP-���N�zH`@1��r"�*_�BX��Q"�/����/����u�,׽��GA-uNF�a�7-��t�bx�s�߂i(=��+jV�xKܝt�x��U�=�����<3�]1B�	�MrA غ7����ډ��3Ns�@&�m)$�V�jՕ�ɻh��T�qX�.\��܆�M(���-�*[�"�V9��|�1�أg��QR�$��hl�YGa]�IԴ�������Կ�/W`������������ɖ�{p���/��N��Һ=+�/)*:�Z,)'0�I��E!��i��~v���}t�l��zXm����ۊ����a�$� �!�ߛ�X�@ӌ]?�����	bN��;�+ĺ�������j���i����r���}�pE�Ƚֳ�;JV>��Vg��VK�y�-�x���[���ɺl�6P�Ij
�o��2�������?4ؼ�y[ѽ�,xYn_؈v
=��ŮW����U����Uk��k.S>X&t�oE~��!N��ȉ�z�f}X�)wZ}c
���ɯ��S�uNݽd�`�֎���+��)ؐ������1��|����i�H^�
�:�:b�1Hpw��|x����_Ҟ@a���Hq�x��m����VC=>f�Pt42�̤(����T�e���fDDϦ��#b��3�	=�-[9<3^J�G=e,�-�΄[�j���� �\�G�Ú`�ӽ��t �m��Z]dH��#w&��(�_7�9{�E̮�}dqzR r!�tߥz��7�3��/w롡T��w�V��e�Y�Iku���W0��G��/�Scu?�Y�'nj#�cN�M�N}�t��Y���Gs� ��U^���b!����U,�jJ{/�=����tW���8�0���:#a�m��I�RW�1�3�\��
�ڏ�"񺇜I��6#���P�V�`�:k�Qt���G��̈́�.���o>6��n;����<݉�_�z"��\_`�e�j��q=�>4lʳ���k?ڠFp@�:��*hԘ[]CGD$�+��vʣe�G�_�f[7�]E9|J���t¥�b�>�bM�W�,ƀ���.\�!����ʐrd���B3L6���nϖ*�E��QŜ��`1_��xÓ۽�wX	Z�m���.�d:��%:�eW���[ �Vdr#�lX��3mK~qOn�L������Qy4�CqDO�����N{�-ȣ�_��=��d{�ǝn�Z�|��`e���H��!@]�� ���/�d�	������"�܃��`ӷj��68%���%k8��#���Cj�W�v�S7��bP�?sJp�z�2��o��#�&��.�`�4�m�T$#��o���*�5�i�
���x9j���"n�<�h)�Py�c�NB9�I��G�J@w��UbP���{)ٽ>� �FЪ�g�c��f��� &~�8�jl����g�I,���#Ďȣ��fBVZ�G����Z	�	���;撀T���Ϗ�*Z�<5��n߾Rs+G+���o��]l� `P�M��-�x6�!*e�� ��0I+�4IA@T�bo@%�^t�㓲��;�t�>ܨ��)���"��hI)�?�ݷ'9���Yu�K
���y��F�$��E&Wy*�t�M�o��R�G�	0lJ:���y�J�:�>Â���`]NB?�T�h��"��Z�3�K�I;*�D�X֖j�{�!�6s!\��y?C1+ycdԭ-S�t^�m�щ�q�3,d��Z����_�ת�B�U�̹�� ^����I�ϰw�O잓���q�Y��s��'�����E�@Ó5��u�d�lq�\�� ��a��\�֭��K(�)"GI<��Mv̔�<�x��#���Vg�".�lע�j8�+ef��N~��H��C���&3\|�0���*h%��9W�ƒ�y�	#�zRZ$�A<�Pn.K��k%yQ�_�֋��ݪL��5�&f`�����l�5������$Z_ٌ���*�@���PY;�"��0�K�^�K���;���tD+��5e9�>�b[_�v3%ۓf:�9����P:��;�u�&bܘ��Uy_�a��Bh?Ǯ20�X�_U�>�HU�!�]qV
m�*�R�i깝�D���'��sf��,�x�/5J�t��&T푧�+��|O�6��B�/{дL�X<.X|�B_[����Jf� ,2�X����4��6#�X��>'�l:�y}09jG�����¿����F�[�����u ��"�B���̩B伭�NjMl5_S�����������E\e�R��\9x�W�U�F�c~|	H��D5<�V�����c4���_@��C��D������a��+tAG"�?l\8�f�ʪ�V�#%=�{����d��u�~����[�R3:�sU��\{`� M,�s�5*e�(�t���1Qh��/Z,��!&�1��C.1}��Ԡ�'^H��ÒXhŚ,�h���jr1��6:"����;�b�	^?�q�y��&s7�>���L U�sx��_ ��fW���G��^���y��e�2��!��~ S��Z��O/���u6��0^��H��x��O{���U4H�^[�H�� ;���f��t.�<�0&a0�M��P�5H�f̷���2�_w���h2�a);�+����C�P�Y�2��L�D�q�Vr�N?���l9������e�R�_�_?�HJvu�����䙹��ڇHOLHk�8Zfσ�������m�5�G.��fd����]�O�	�#Ĵ�?)��d���>+i1��Q6�������Yhh�I��y���bx�0�a�����VQ���m����P�4?|`� �:-B�� ��׍m�g�-�%צ���$�7�|\��mWA�m���c���,�tL[��w�݊�~&�}f����ێa�/�Sߢ�����B���ɋJ�nhf�`|f���m7�At��Wס u�����y�%�qV4܏�������D��v]��x�������ٯ�^Q9T�d!d8���<R���B2t�P +�V��Ȼ����q�1�fX�����VF��&�t�����OOψN��W ,NY��Y���N'Id���`��ۣ�y��b��l�{\y{I�S VU)II�xl�&��p����|!;�B�=��7aS�gK���׽�Ff���^F��&Ԥ$����d���Fb7f��;�f�9��Gr�Mh#��ڣ#�4���>?2,δ@gNX���i!=�Y\�QzEA�u�$��ͅ
-G$����Қ��F��;��I���#����?���o1��^x����R��|����G��Na�(f��+Űj�|�~�����&�[ƘZ�*��$X$�UmP+3�G���w�-s�&o�E�Ti�AgHbḚ�ۏ1z�Ipd�����e����3!�%_�?�4~M�,?nx&��6{�$-�S���еȂ��-L�]_p��{ؼ��e+�!E^�j)��m$.��^��n�]���e6�=���#� �3���2�H%!5cv2�攝5F<
5Q����:�4�~D�լ%�G%Q����ծ����/�gД����t�B3wqGJ�"pd/�}ܓ�����J�GWgy��!��Ȃ�������`�Q�ձ!�?.b݋,�z�2 ;�����C�Ì8D��l7�H���R�-�O=��	�X^���K�Ł��`8�ѡ~���Z�-ƈ8[���#2a��x��kG��������%K%(��.U�~ve>�k��@��� �>Y�����o�iCq䘊�:w����\A���N�X�En=��PS4��v�� �����XQ�Wx�rhеM*17��0�i\���)yXHe����Πɥ�Yfi�+�-��"&Ccl^�[�V�LV�+U<8e�#�h�7د%�9�O�T��{/���:�^��A�VU-0���`S uy3����S�iO2�{���M��ϚS�� ��#9s���lOy������!�����JGt��ŵ�f��T'�CH�O�@D��h��J{���@��x&\С���uk��hy�}W(��eM)e@_�{����Wq�G��tS��|5P�� �m!�Ø��ZR	��	t��a̅�ŉ�q-�a}A�f�x�#{P�F�mi]�C�������)�R��W.y��rFH�g�tp���o5x�s�y��M��4l����h��ɗ����1\؄��ȵ�`���	cM�첦^!^�z��u�C4��/˅{�H�YG�^�vu���\��_���<��0k�W�jFS�!�LW���<��,S�H��w���J�~���w�$`2�y�4���7�1����� �i w2��EL�i���0�!9���c�vj]"����?]2��F�b�c�F;��5bք�ɟ԰Ni�-�d���<w W
��%=nh��X]C���ŜFQ�Dʀ˗��SB�,��o��j�;.(���q��p;�	@�D($������5~��?����=���K�p�C���]X�.������6N7�R����R�z^�C�x2�]
�(�����_e��a�-y&U,�7:�20l�H$�#�[��I0W	�l>DG�X�u���"�A�tf�#�(A�lҼ�B�D
C��X�cb$�L"x��t��.�5���Hr��z�ʰ�k��\r�1�XΩ��� �����zz ������q(�ݗr��	��g vg�����}��y�룈��Qs	+t���l�ޱw��J�z��Ђ��Y���\�~QL���Ŝ������~:I8- Lu��.<,�;�O���b]}���kz�=������vó������%�����Y_�h��W´�d��B�y�l y���.�_=u�Fa�`A��������ʅ�) �W����HH�b��9�HY��
�&�O����꣟���c�M���Gy�߰�k�r�Lʢ�k�`�a���ҥNlqN��e����\�.&�ԯ�����֕~*��+�ܞ���h\0^r�}�!EՊHj%��M��{��x��Y����3d��B��dٜ�v9�0v��P�0�;�A#ڸ/���C5�哕>���A��*����[�FZ����@:ik����#u��qw >�29�����4b�,L��n��YSu�E�n)w@��N������o�hwD�@�7&�[�OPCXS�ԆC}E/�����/�����u�)J/�� י�]*��S��lq��@ި�w�#<[� m,}a�ǴԎ���FL�\K��pO��\&��!�u���tz�@!���鶌U��BeoD��UI9������NBS�%��`R/�i���S�\N���Y	��B�Ŵ�3�z�#M8��X���&����2K5�j�<]v��ݥ������-���θ�*����0�}�Z�f���!�;76�l(N��7y��;���؍�2�g� :�0,��}`�ƌҢ������M%��<�0���79ÐC�1�!�����MTh\0��Ѩ+�J����0�20�A��+h��uIy��Li��4h�<e�7t�B�n���掃�*��p��ŀ��;��ٜ���5`�A/��/�ԥL`[���Z�{��Pz$(�P��v��4qLyn��[�m�7�aֱ������Λ��B@�⌥Ng��o�*Ъ����kç����'p�U�$�1���̹E'ä�.c�Q�*Z���Ad�������(���L�'�(��OW����\0G��N�1EL��ܕ�Q'镁9��b8�F[��Tl�y7����m�k�(�,p4���%@t���۷A��+�cD����r��:e^�TH�d�ycڄ�8�E���=ش�t��B�󌉎�����Խu�y2c2o�o3���{&"�@�'S�)Q3)�g��n���#Šޕ��o/|�V�A��P�;�j��b���Ng��t��C�_�E�1��c�F�]�
ɀ���W����W�����J֞XQ ��d�o�)߫m�uɕ��,�l�z�I9�X�D{˷�$=�6����䈷�nFڪ]�6���b�m
��~;��R��	���w=}˲M��K/��Xe>p�{��>�x����
$Y?JQC�WD�yV{>A�䫘�q�=:2���jQHUk}�X��؅lHP�O@���T}�}��T��DL��3VQ����@���B8l��n�X������r�J���bF����v"1�V:��y& �Dq�f�u������ �e���J��қ�u���q#4�����o.򨽫�.V#u���K�T��<T^���:�Y�٨z)��%�X�vu�� �@���LǴ^D�mٟ�1̠�+P2ԦY@�qKaH�8�a�.�8Ύ2��R(Eu�I�] ��'�Td�a��KFD�2���O�+�щ3�	>~�;�����M+�������BX�3E:�=04Ymh�
�f��t�o��)_��R���a�1�&ʷn�PӒ���v�\��t��0�,G�@�ό�j{��Ş��LLX�Nj���A8�����5�3Lkm�{,/�۷#��Z��2�	��N��