��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t�������.NT�ɯQ�_�EY�����]|�=�Ăt��@��{D;ӸBr���J��;��?�͠�j\i�ş%m&j��?v�W���tF��NO1���?!T�Tg�U-�(�	Z1�B�#q�@�;<t��:�[-���&��5/(���{���i�9�о=�%}�~BW.p~+`�l�`�Y#<y�{ˢ�0GS6�����P,�pʄ������9�5� 0�X��ª@���>DS_���6�Y��?�T��V ���4�$X�__�w߅Qo�;�g)?�Z��Ʈ$D�V�{\S`�&����ܜ��OYo]�9���$RH˰�;G�&k�<��,_�t$)�2,i�z8�8����I[3.����sϋd37���թ�Us���ѱ([^�/�9�V`��չ ��N�󸁧:�y9v�q��2��a U���(�s��i��o���:jal�b���3 ����_
X�)Dۅ:����JV��Yd���p��"��\�h�
�&�eT�mZ��j{�%��u�Ig�ҳ�)Md�[њ�2K�8��ꈃ@��G9��h�ۆ�ɖ��$C�����J�O3)2/7�-�z��)먀?�_�V�1�\y�̶$ȓ���sX<��Ym˙Lq�Ry�1S��,��S��`ۊ��� 뢖��_t=Mg[��T�M�<l'M�nZ���؃��C����|�0Xy�s���p��ZJ���\�Uh@�T@1�/D�f����|�|�}�sѼPM`긻7 H�@���4���2՚����C�M
0�H���� JW�tNP�C��0���V����$�0��R��kՐ`�G��w�Au�ƹF~F��+Vs������&s�j8Z�l��	1?��˽�Za� `��.�_(BL���"���%�R�R��)�f����(C 
]����N�7]��Nyw���"� �����?�;ok*�����,�o*͡
:[G���b.�0�|>ja��F>�.�����N0��ٶެ�V�w�Q
������Ҵ� �y��z	-/�y�C��ہq���0���{:q\km���)4�^Nچ���U������g`�&����M����{�J�Fm�dC)�b�MH�8��p�eP��a��!Z��I������e�����u�CE�����>� ��W8H�o�?�}��jO=���NI;���zE2�d�x�s�b[�?��[�F����F4᪠��:Ne���@��<�ƿ�t\��3�M5����Q��7��{� ք
�lv��eǂ`����ŕ�?��^REF��TjK~��0f�V,�����у�2^��*�D*�~��3p'`�����C_��\���>A|o����bC�it©�/�Ft���6�1��+��ffl�a���$u�x�{'	D!�܌�	:�j���g�P�����P�Z��
 N^�� =N
�d@-95~���rb�t]^�*s,үz=���?��3{�5��k0����y�2���&�%�77�6�I���y����]���a#c�iv�\_"��(A��LM~	�n���p}fw�pQ�"u��-��#j���*n�C�\rS"�?����{9�a�?]����?�-E�0ߨ"��(�������{�-	�>����Q�"a�O(��c���T�C;��[��o�����~�l�����y/�¢ϭ�K�r�M��1�ױ�y�vF"��B?)�C�*�ex�e~�W��qf��L�#_g�8=y�����L���f|�m�<���5?�^��o�?Dl�6���z���{�L���2P����k�46��ոN��g*n,yUqlk���!
#*rW�s�A�U��Z��Jس��4rz�EΝY���r���B��Ђ��&	j�?c>î+ qh�3��pd�/=����V�R0�	����K[�ʯ(^�S�H��'�\�����m2|?ᔎW�ڵ<�p{��h��-���D�s����q�$n�5½% α���J�	/��x�"�M���ٖ����z�b�k	��dۖF!�7L�{��e��<�Tw�1[�&<0ť��ˤcv����='؆��+`t�������)�r�ESXsf�FP��w`����PT���4.,�L����h�Y��u5��eY7kʹĥ����2��qH�h�,��zvv�UBS���b�m>}��S�fB�)�h)�u�Z�G0��ZzB67�P���&��>�W�c=ޠ��?ۅPs9i6�'�Uu��ʻ �d:� @zƧ��(���߃Up%�����(ՇNX��´Y���4�m�鶦��骾��|T�ڀH��	M���'�F�^zL���C�O	�-���J�d��w\�ر׮X締`8�A��4�h�R���q�Bq�Y���6;���4�˷ww��qEU۩�+�Te�*E�P�3p��'��eb�K5��5'!	�����oʳ~�G$��JW�%HM7]C�˦�e`�Ō��m�m�����W��G���w�R��6zSJ���q>r�����xәNuΦY������6�0D����"��]�P�>�ۆ����J�0�4E�7__E�Xp"�]UB�΢����캦T�t�/��`X��.f̆�`���4�޳�ٜ�'���L�:����P?��MЎ:UBl��>;�ww���C���d��j���]�mϖ
Q=�a�X$��x[�G���^L�v�%g�e�Nɇ=��iS�K.ހ��*��D4�?�ܚ`h���%���y&5h~�=�y�[��QM@����K����B�sl�ę�L������h�;����1!��QҴ�%���*ү�Cˆ%"��´済��L���Kz�HoVg{G߇�b�d'�a�H��c���j����xW|�??�5��~T��崲X~zu��$��=���6K��O	��I�B��ܣ��������3ǵkI�����T�wP��G��`�9��ǖ�h�����ډ��Kb�/����đ��V�5�X�&)IS�Gr���珞�^<"�����]v{�h�6ߛ	-��m*gyS�1y@���{���4Rѱ�(�m!y�y�H7�ua���R#W�����ϋ��8Nw?��B��/��^av|��|�
�	X +��&וS��V���Ŷ��&7��7��L�@��ՑZw��c>5�w��k-�k'�X��֭���	�b���������Ǟ�:������]t:�;߆v�(۳���?�W�t��v��@@�(�Y�Q0h������l޽!|=mҏ!��"G����o)�29�n�h�C��"�&��0 	��]KAh!�or��i�s3X���&ʺ�����Js��~�M�KEuc�������<6GԒf�}xܨ�42P�� ��1�M+�bL`1�d�*��tK��uR[m����}/�=�Gߚ~yG=kr����+<���R~l��G��U�(G{fhL^(��FCn�R賮�)���J�z�9L�����i"ɔ�'�Γh����V'�РO�aߨ�R'�l�0̴o��2wW9�Mh�38������I���� �	_�Jv���;)��b�{0�J?��܌i&�����`���?�+��u([8į�N"�;�����+���d����D�^/�m���&�R�g�.ѲO��1�.�/�]>pL��j�h����n�Z�$B�p��I�@qJ0�Pb*Bv���j�%��c���@C���i|�%���j,�y���� ���6.b9���O�ޚTu���F��~F�a��,����D����C��6%�̽Z�؃ ��1�m�S5(�dco�,�Xn%���T�/J�zm则^;�[n��M�����ԋ��̤T�e�*@��KaP��Vr#�
	x1z��u�|�{ƣHNA��"E3t�%JP��)8*s��#�p�Ch/u��|�-�-�f�B?˅_��Nq�m��Е|�KLh���R�Aȓ�U�k�5��*H~Չ�^ض��e0%��"�}!�9U��.~�o�E����t��][��W�ô�����%ؚ��Y`�S0zl��:=�8<�����u��:}�&�
������,������xR��og�!(�^��j�o�Yͅ��N�h-o��~�8c�u�gh�+��<��%�ѐ1��V��q�'�S?������v� �?�١b_(]s=[W��:|�vA����>`��:�GMJ^8����Z~RVi�����x�H��e@����������,�I���F�\rp&Zb���G0����]���b�`z-_/w�^5�X���ՋHɦW�l@64&I��)X�1�L1�<D����c���� M�s�V�~�	�V��,���wȣ�w���U^����,;ъ� o�SD�K<�-���{���)����#pY�_�.��Q��2�5~�g�<<���G�@u`���P'���y���U�U_xM�����ѢOpO�%JO�i��I���`�G:�Fm�̺[��>&��� z��1���c��1A��h�O^� yDv���eG����z�$�]�>���q�d?�x�`b�KHz�Jl":_�M�j�LgJ@��H-�0�r(���?uYo`�7?Q�Hu%ô�ƯaQx�a5ћ�D:���m�Z@�.Iسٯ8�÷��r��J�+��*G�&�B·��V�t�y�z;'��;&��R_{j�.�`�F�x��~��� �s��ީ�	>F�]H�X�	za���.�Y��К�Sn����ĀVF��+0�ʖFN5i_�7�։j�p��yZ`�S��1{A�R�@AB�x/�!m�k���B8;�B���g"-�B<�豭���ƭc��Hs��JS�o��!�U�O��m�Н�2v�5s�Wx
q�	'ěY���t�r%�`��\�֣�&6��(�	x6{m���"� ��(�͘��i\��n��d� �tQ�2	e������0���[�#����N��gn��S�X�a��=�vs�<�Wq�<�_]F{���&�Tu%�D��W�i\�t�K7��j�� iig �tx� z��B���f����Q{=���=Z連���W�����	ӊ��i�:�6t)_���u+��_ 5 ,w�8xe�d$ �t(u�c�!8��`��d/R�v(���e����;	N\D��T�û Ҡ{f���,o��+ׅ@�:m�Zr	�.ѣ�29�C���`k�F������tB�Z��i@1ò��Q���A���rW���-!�`�kr��vISӌo�݊�����o��a U���`�i����-�% u��n��S`�B����Y^����m��@���ҔNY�O"*�ܹ��̗Z�3��n�Ґ�F�n�����}9T� ��{�՜#�$m��Om)s�r����#����M���sF ����>�d��ݓ%n��pP�c��eN֥�����b�T�؊#%��1d�[�)#����|�Kk���վ��D��WF��Ī���8�ܾǎ�=�S4�?���\a�}Y�M2�]������,���S�Ck�B����Y�Y��pU5���,yl�����X�̆Y�H��̰S���O'Jbr�:�@�|.�i�O�@�t���1��6����� ���׼��s�Z
��}JOIf](�>Ӡx}@ڗQ{�&J��s0��c�^�F���e��G��4u�˲5�'~�!�R�Y�$�K��>����X�d#$�sU'6ґC|f��X��N��(i�w�oOx�%���!ĜDl��墕|�{�g�Rs.��R��5w�?���L�N�xf
�j �G����ͺ����BD�u���K};(��|��ҜsY��z׺��l](���~�x����Bs�<u�'�\V9Z+m*;�[pҹ��L�y�d	�5�P�m7Y�ʐ��S�~F�av��y�\�G���3�oY�p�
����xh?����|z��>��P�+z.��"}h�ƣ�~���44op ��i�/Y�۬h��㒟}WT��?V���
L��D�%���[�`�I��Yϵ�LFA\��=6VK�:�߾<���տ��ߥ3�N�%�i%�M�A��N�{�]o]M�� �����.ȅ�Gby-�w!�A��5�@o�i�n�u�Z��#����H�{�']�ȼ�2i����2qW�AkT�@����^F���j���IgfN<�����N���P��{�:l�@T@������c�<��Țbt`��ok��R��%����UB;��#��s���_]���}�WN��F _(c���Q���N�M����V!2g�����V��5��� ���yg,�[BY�R�LM_���Q���! W�BZ�`U��N;��I�!C<�KT�����!g^�,6}��p��s�<���&F4�9���6[<d(@�������Nwx����oXqWp2͎�
�n�x�N�W�2�|�r��eڊtKyO����G>ԡ�7a2�ߍ#�he4�mI���m�qJ����9���I��~W!ɛEMH��@��YB��7�}�V�qaV
�!��F��q�"��t�����ƁB�%�%��U�lv�P�D�s�������_7=���c2����݈R�Ņk�b��Ϛ�H
A$JRu���gw�����,����U.E��V�F�=�Ш�ۭ&O��$�DQ�|H��Iq�0�!1�6�c���d��R�P���|�O�h�b������#�vN`����R��G��b�xRoa�Z��q&��V?�A�ò\Ҳ{&)��VA�rkt�?+E~�}ću�_��b�0RH�A�ނ���xX�4t���f5���!�R{1O���.(p�>mԆ�}}%Z[�]�����߷�h��?�<���^��r%s������� &���V��5��w��Ƌ��,�А�t/�ΉYtY2����C�T����K�yW?$�SI1��4�-��b�l�G,�hwmŰ��{J`������p��`��;�~ӟ�G�YTd)LѾZ7�{$����U���Hi(D;�5�.�k)���SB My�[r�1�RF'z(֜0�I�<�d��>J��5��X�8]9�w�0����̴�x���{������T���t�{���2E����n�@X�Rx�5��4ą�% ��t�:�VЫY���~��[~� ˧$o\	h��~9��.�b�,#e�mz�H�
n�1�R<�E���%T��LIЛ;+ۊjX�B�1V�h=g���n�[�>��>~�����
��̣�2���'�T�3�0'�&�p��g�ޙ ��-�q��L��#�|V*R��5>�*Q����ň�ʼ��L�ۡ�D����#��Q�=�����H ���6d�Ň?�"ђ��:f=:�Lm�v��3y��w���DU�M6���y6e=�떳��%Y�ʽ�>������(�E�u�g_O��X�^_,�f����p������M�!+�e�)X�}�j0� �3�P���hG���*��X��@�o�O�F��`�v鳔RG�/�ɓ�59�}S}=�]J��d�� fC[��G?�FѤf6� I�Pj�_Ü9���R��%������^��Pl���Ҩ�r�oOb^%r��S�ۧ��ke�!���_�XI�����;1�w�bކ����z	-LK�������qU��O�!fҝ#U���,�>���\������W#]p~Ԟ��˔�EȪMy�H�H�@�_�Zj�]-�~b9���4���6�>	�Q�Uqv(|:��~��C�T;��������GZLlPcL�:��]h��5n�lp�Q��؈�w*���^��	8Aa�ɤ@����ā�fȜ#�����FSڏ9B��[��OZ��joSH�,���]L�"��.�Ԓ�ƨɉ,��pԗ��d'��_���1��C>�搩CЩ ��$g�.��M��N�,��ܢS������)q5 
�V��s��J��s���$ku9�,�AB,C3�6f.O*��N�7�(؀ѯkU_��Z��2vT=�&D/-��jƟ��5ۿ'�?W�Q,5��X��"�.����.����ڨRŌ��`K�3�^���Y�����uΎl�zf(X_"�pAK=�؂8��yŖE�h;�N^�˧�?���h�;m1��"�SύǭR�!���րS>T��#$;ong�C�����*�g�1���t��X_:5r�5Yy������m�6�K�̥V�8M��b��4��\l��4Y�"xJ�D�KbV�=�q]C��c��'�Ԥ+���]�Mef�����}�e͐��q��_aVg����	���JRV.�W�_5���"jX�nr�/�����ӡ�n#"�;�?�B���cJ7���(3\,�hY�ؘ��\'���)�������rJ�-�<�^��q��0�~�Frk�ǂd���F�98���`���fR�x�]��ߖׇe��k�zs=�k�2ph�KC+���=U�q��$�ϥjW��w%4�R����B� !����~`I�B�쪁����.d���)=��E��s�rq�T���K�k_��Y�f��bg3�>��s�橓_+�J\�z�<Hq��+>���tAyuK�1з4e�{�}N�|T�o�%Y�\���0����(l�Y�$f��?�2�
�Xf(��9�kD�{����C��葜KqZ��.�*���p�"B(�� l�4���E�6t����!�v<���)�����q<DB��Q��o[�.琣쨑?J���f���d?�ыD���t���(���ԥ�WK��w���/&9�
E�U>��}��	J�~�0\-Oo"��l1��5�#��A�p0�ziP���M���:#ќ�_�^�QN����>��/?"��E*�CN�k��l��Z�+�+s�)����^h�Ͼe�W�Y��%A)�RAs���|G~�+SΝ�g��,�#V�Ҽd����݌�5X=�� Q�*�x.��a��F��v�UP͵��s�8��ov�M��'