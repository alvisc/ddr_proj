��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t�������.NT�ɯQ�_�EY�����]|�=�Ăt��@��{D;ӸBr���J��;��?�͠�j\i�ş%m&j��?v�W���tF��NO1���?!T�Tg�U-�(�	Z1��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC. �,"��'��g�	���:)J�U��>F���\(V��S�Y0�$�Sv�ջ'�c�@��mt+�:4�.�Y��X\
��z*WR�||"�i"�����ᓇ!�I+��_�Ph�5�5&ig @���bl����4Lꭱ�jy1Q7�r\X3p �Y|���u	��[e�Ƕ����+Ƴ�K��$[{��ha
����6�{/c�wD��J��R, `�s�K�7W �fr�!o��;b���A�ͺ� ����\��o�XŖ��N+�}j%j��O~m!�׹еv��>�r�6������v�� y,ۆ�]@}�:�e��=���I� �~��czK�PB��H���z8H6��7R_&�2�m�Z�tܷQ�2%��C�Hf '׃O_ځa,�ؤ�<3~.;|J�R	�j�*���)�4Rkh�����J���� ��B�6�7QWU��>B��;�cF�2�n�L�c��8�0�;��Ů9��k�|��Tm��J�iԬ�T��D�l�uC0-�Q2Ұ�ܸ�3(���t0��Id$�L�-�Gb�	kj��D��`�U׮�Pw�X�.������2����(�䧀���-E}˯�8p�nQ��?\��nU�N�����u���s��y��@�r�-���4s M���%8�u���'%'d���,K��b��K�s�Ьw���r=�45��C�:�%� ;Cm���q�����Q�闰�^�@3p�I4�4��M�a��ڿ$�;�c�Us�
��Vf������xV�~�W񴔋C�3�ɢ?�y{�a�#B�`Gd�e��Ƙ�gX��{�<�*}�������?t��`^�t���2�)H
 �v*(��II�uAƚ%�R�(_O:���k�hg� ��7����&w�<Ső�B@��x��ȷ���=!e\�5��<ۻn���a��2* ^��fy���ش�n����M�_�l*���S�hpA5z����m�g��%��I[ZI��R�xqe[�8LSêM���7[�>��%�T�z�?� M'&�?���:�E]$-�J��-����%�,���?bK^ ��)Lw1Anq����<Y iu��,���%~�NL�w�G��0-e�@��\�^Z��):K����$`b��O��H8�i"�	�7+���0����zJˏO��cߕ�_#Ok������v����>�E��G����'m^�Z�,
B����u4���)2H'���Vw�v!���T0�ϕ0O��w���Yp-
%�^����Fv8Kt���ꞌ�2�ј������N҅Rggް��,�a�Hw!ﱳ����F���?	y���>�޼�n���f8|]p�8�*B�����|�	m�����')/7�G�y��u>������|eJ���T˙8:dг�s��P �(U>�A�Ө3��ۉ�3�2Vb�?��T��9�/�n�(+k�		5'���M�H���X��l/��V�vOi
���1Mn�-���k �mk@o�p&U�����x�z��V����4���9�|Þ�����bln@��>��6$s�1��9/�͍״�(?S�"F��A
�D�]���9�ș�Y��0��QD��O����;����7	@9.T�P�Lj1)$���DA���4��������'&
Ɛx���+�S�4@��W�6��֞W��m�b�a�Hi�G�
�=ܴf�o��U�(Z��Ǿ@���h�)��!,,�(a�rHV��h��2;�n�f���
�z�ۥ,���%�n��ŎI<�0��2+};��\g��9*��^[J;n��l���,X�e�p��5)��í�<�\Q´w��>���[�{��i���PJ&�)ni�PbN���7��g	<��HR���Ҹy}�T����J�;y�3�Sja�w�(lM>.#�g�E�Գ�����1m?#�
�1o+2
�,3��r	k!:��E��6~!.F���1�T�<��|�!XƖI�()9҆�l����T�f!�	~JLd/�I��[f�)�W0��`͔I�}/��.���zW���n�Eg�s<�<|��
I�&`�T�jo�7��D1�7x%|j��@߰XI��4�ʼ'5�5�M�@�j�
vV� ��Fr0�'���,3G���W8"�03
��8xI�7�]��uR���g�u!NT�њ�SL�1q|S��	��n���1�+�=�2��~�K�X��IA*���?W��~HL�:h�U�K�9��F��9:r��k�)�o̟k�T����V�((���p*0����2���_	L��|s?�etK}P6Da�=*�P��V�+�]V׈�b�;b�m���r��%/�����3L���l�a�)��N~n�(��#-40�d��L�KS"֏��<�[i���,g�A�=�ܐ��;�$����o���iQ��Đ�ڙ����A��,�I�2>��)0���z}�G���[#s��ro�.����~����p�
TS�?�Ŕ����_�I)k	N5P�'y^����g<o=r�\��7��K�3�Г{�4s����2y���U�ZA�����3�D����,����2�_iga���X��s��c�T��O�qG>��W�m��) Q3(be��izw�Kx�==a{�?������8�p���b�y^�&�E�O��n���)�GJL�R�X���P"���� }^�\�8�%f䮛�x�`� Y\�̦���%�vf�����EWOCЪ	Pէ�~�����Dt����-�l	A*ʽ5��ں�~�^�w�la���h�(4�������杈��W<a}���GL�oK��t�N���4��w=���	��QS?��p�F%~g��I'����om�XZ�&!������>"�aP�mL�l�n���n���Uf���e_d��J8͋�Z_C
"�5(0���O�{S>];O?q�s��c}E�&���4Ly��\BJ��<;�ӪΊF� >����Hoj�����~�����u���LK�M#����NF�]&/xj�����%t��g�U���q����J�] 8��:lM��t�k�2����Nn'�1�;U`ئ��ӏ~����������<���-�R�챌�2#�:��K���]ظ~��1W��+%�eY.�S�z_K�|_<�8���`�(���^��[ߟ�09�$<��k�a>��j��lE	�w�"��_	�/���>c�!1�f����8�䝉Fj6�"�.�cY0�m���f`U�ehd���h'��a�1�ŻM�葄�u�Z�ɩ�$� �a���H�0���F(��a�,�/�_L4�#x���"܇�l+T��ӥ��)g����4>'�q�'EB�@�502z�K�d�0!�m�欭�!}l�Ъ$3�'ES�F����1�O�D��u�L�W��|�Tr)zuq�(��B����U�|������+�>��B��"���twuO�+쟲Xw�sf~}���3��l��G�oZ��r!������)�6 &�����%�-��(P��H�/kɸ���x��
#I�[~���t�1:P�\�׎�ǔX4��[�ce����D7aʒlZ�i��)�Rkg+԰�R/č@��KWyB��N�����	�4�w���{RY;r���#�!����Q�%�9�V��D���?�ݩUQ{��#��mn-�C,,.�9j�W�߫Xp�_��C�&��[	>�ǁ��$F�f�I,/::#�H����ԍ��y���ѩx~�HO����{ҟ>�*q?X��4��x�K�m�i��������Ih������3��SEǂ]�K���9������ �ˌ]�Ң>�A��KS��/ģ0e`�:lH�KT{��`^��5�
7�ːJ�w�f��a���N1^�-����f���U����[ ����L0E&�c����a��/�7��➽]��ڒ�ӌ�E#�[5Y���V����np�}�2b�p�2�h�A���'��=�Ѫ뵮�}��1\�y*��T�+�V�b�Iӑ�"�|%�F_7K��f��s�rCF�a��@G���.�������1*�`�NqJ����X���(����ǃ���`�bp�
C�ێ�VMn`���2'�3w��j
7���6��.�
Y+�r/ՄS�;8���߫L�Ŏ� n)N�_d�?x��J��Y}]���#��0��L�l-�qb�Ϊߡ�+�&6�΍f΋�chOZ��u��ʂ�8�6H���[l����� ��1�Z�o��Gs�k�H^U6�i�Y���p�t�9�ð�4t�]�r�Ƿx6C#�i�1a���ُ:-�e�<����GM�O�5�����~�aԵ��j�_�@�A��Zz�f[�yB���/��k�m��+F���Z����{��&47?J~:�qWt^�ꙻNu���"O���({̺m=T��������Hep��[ C��2p���ET(�����M���̮k�5q�gܟ���9�S����m�����s����+��>�b'"E:�y�R�W�@^~�
�2p�R5K:�o�'A�?$�?]�:�~�门y���9�1�g�u��-â���_���(�H�H���(�T��s�M,����T̄��ōB�8/O���\���٥q�a#��1��x�.��Ō��0����S1�b ��W�jM'��Fu�m%��-�٫u�]�x/󨈪6�F�k�@	1* �'U4��8[�����yO����B��@_���h����ͧ��,�C�>x�H�<Y;�O�:�٫]b
�6be��?�կ�0>�.���P=�VU$%H=���RC[����
�_�V3�}b�����h���'uw�;G˦�����ܔ�8
�t��a��S1}t��
�~,��Y� "�����J��M��O�sŶ����7�3��P��9�+�ڲ������Vm{���&|��밭H�(�3x3��Fe�Gd1�aD�z�ZjpJ�6�~M̡&�G#a�&!O>8w�sz�^o架e�@����,�Vm$x��+�r���*[��yK闋r�$l��tPZ�P������C�����'��6殑�r�N���*�9t݌��}�}7`o�]N|�"����D�Q���e�'��;};���_뢅�AMϊ7��k����v�z�I�Y��$��Gd�?�2gXH��A����o0u�ˆ�m�ati�<ff��
������T�U�ҏ'�YF)�n���X|�p�$��~m��aE���U�1H���߀�N��l@nf��g