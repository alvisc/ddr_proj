��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t�������.NT�ɯQ�_�EY�����]|�=�Ăt��@��{D;ӸBr���J��;��?�͠�j\i�ş%m&j��?v�W���tF��NO1���?!T�Tg�U-�(�	Z1��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC. �,"��'��g�	���:)J�U��>F���\(V��S�Y0�$�Sv�ջ'�c�@��mt+�:4�.�Y��X\
��z*WR�||"�i"�����ᓇ!�I+��_�Ph�5�5&ig @���bl����4Lꭱ�jy1Q7�r\X3p �Y|���u	��[e�Ƕ����+Ƴ�K��$[{��ha
����6�{/c�wD��J��R, `�s�K�ų��/���_�^�r6}F���XTcFǲ�r�t[e7l^�Eu�n�=�"X�崺%����ή�6V$4���,-O��0:��(5���]������[��/1��-�F�	G�ಥ�}��၈��`�s�smyo��9��5�ܧ6�(1E��
�����ɸ�Bo�Uޣ���]�9���hg���̌��<�(��A[r���7~�C%��F��d�0��e�
p.�Y�UD�9��!��!�堕�be��~�X�}6�4�	3�f�Ć��E�|�f���O׈	J�<�	g'ǩ <.�b���rR���׏6���'�b ��t7��Y�<5�V�|̮`��\�k?����B`3��*Ϳ��q�{0�8Q+�`��{Ą���Nѯ*��X)it؝��qJB{����4���mV���vU3l,+[*�=��>�\G����`�J�&� +�چ�4���Z�`/��g�3E����6o�n1���������-�z���FxD�Ҏ���ߍ8�'V����,�� Ϫ�&��!����ړO�#��`Z2�m�@�ͨ>?P�q��Im��U7Y�w����
<�B�3��O�*�L��+�J�O�"*Wj���I)�	wF�B����k@�Ӡ�Q��'��T``t�������a�u���xLW�f�Eu>h"�s|Y�4�=�+I���0���h炒�3v�(���N4"&�V�����~�e�I�'x�z5U�d��K�+���K=
Wׅ����y���F;����̂�}RZ�{%����ޔ�K�y��nϵ�ebX'���:ǵ;��"��iw��K�q
��ƋϬo��������a�E`�!�Ο� ��r5OG�����ڎ��z��H���+���~�D�+S��_�5W���R2G{dWf1�+��\��]�;,-�ɕ6�|��&(yW�&�쥓��l���D]�"��H��K���" k��h�a��2�(�u�����h��>��|�������p͚/�v5���H�����6�6\�,�Mo�i-y}��K[͜�G2OU��~<{�������$�c_�ݻE����Ձ�`���d�\��CNp��rs������M�u���O.����?H(�M�'ݔ�	�4چ�煉##DΉd���y{�KjE��ʋi1Gg�����hq=��c����W7גs�r=ǋq��	����E�>5�O�6:(T��پ$T���6�Q�{݀zu���1��샒Ш�E���F���T�3K��i��&�QZ�/��4s�f���=��g�C�����'��$��LB��v���(Pښ�3r��z�����h�?j̰MɊ	�H^�W�b	��s=S��Sz�9s�X�/��y��i��o��.���pJ�C�n�ج'�� �'p\�(;�F��m��d��Ѡ��ck���"������Xȷc��<&�ڮ8�}'m@/	� 43O?B������E��웩��B�8�n�D	y;�ޅt[�7�Uٍxs�9�� 7�Hծ�&�~m����E�`��~8�'�݁��*���Ue����b��S��bd��`e8�!Y�� Ԧʬ,R"�\����\7ml��Z�"d�*<�ƛ�T�y���H�抺������X/�GD��P��A��h!ٹ8�u��<������v���'\�k�l�i��u���1А@�N���`��κ��&��Ā����غv~m���Q� ��Cck��9~�^�o��Y�|�������t2�f���7�Դ��_.�!G��ԭ]���j�$��az��NJ.����4'�4�a�[�iW�c폍I��Y����I��'y�]�@�V�Т�@�(�Khff���E[g�4&�l�ӥ�I+�,Ѝ���Hg�������,�r]����\!:�rds���̶[Z]����9�ѯ4( 1
�o�s}å��ã�m�TI�^�8*i�QsA�x ���?�*�?U߭�ˎ��֏��{I�5e� �,ɓi�}lb*�G��*�>Y���.>픋ʘ��L�.<P_Q���DIJ�I3��R巶=���^�S���gړ{4%]��&�o��]떷�!>�S��"���i�N���+�6N��k��rp�h�����n�~�rc�ք���D.�׈��\��)Km�Al	�n̔ה_�	����Yl�ub��!�I�3��eL�q�7X2��.�b���5�$�2K�9�6Д������tQX��y�%Zb�|3Tȷ���Ң�	�̖\̾��\N�43�yW#��j�c*U�ř(ڠ�L�_B��9�U����'T ]�3sP��-D��m�Y�.�u���Hc��g/�fUY���&��cÄ�Z�JW��ؕw�$��GZ����bs�N��Ս��������6|X�>���Ǿ�^�8��t��*hh<E�S7%F��}��)� )�6��u�LS��шw#"k�$��Y��H*"Pߒ��V��E�͠V5�(���&��
����-܀)�����'�=�h"�H�.��Y��U}�&�Od�+Tʼ@�~�����5Tc
n>�,3V��B��T�C��T�P�G�|sQ~z��J����s�5�� <%��<�稍+nS����I�_��!�(��IZ����4��I��|��{�f_�V3P���o�n^��R�����N${#�{2�cl��/MV˒Wl+��VoGM��5,�Z@Hc0�VB(��걨M���1��&LF��;�A��"�OzRy�G/��j�� G�`R�L,[��������h�Ecn��\"b0�R�¡�8d����䊡�=�����"Ъꋺn���wNy��~k$MR�~�v�1@�}����JK0���:d?ڸ�nTK��#���U��*e��W��z="�d����+���S{�E�5��)� `o����k"�).���!N˃Y�Q(3��%t+F�і����k�-K����^��t�b�(��p{Ŝ�9��%˧����/��$������UF�����&���7(�Qᔒ����)mz���!� �PDЩ"��������k�����:PdP���V����>���/�8(��Z`��%Đ�7fQ�M�U�	�=�����X�o�E�^`���F�Ny�=�a�����8�B��§�����Fu�w�
,�yܨ:���k